//
// File: hvl_axi4_2x2_fabric_qvip.sv
//
// Generated from Mentor VIP Configurator (20160818)
// Generated using Mentor VIP Library ( 10_5b : 09/04/2016:09:24 )
//
module hvl_axi4_2x2_fabric_qvip;
    import uvm_pkg::*;
    
    `include "test_packages.svh"
    
    initial
    begin
        run_test();
    end

endmodule: hvl_axi4_2x2_fabric_qvip
