//
// File: test_packages.svh
//
// Generated from Mentor VIP Configurator (20200402)
// Generated using Mentor VIP Library ( 2020.2 : 04/19/2020:18:58 )
//

import qvip_agents_test_pkg::*;

// Add other packages here as required
