    Mac OS X            	   2   �      �                                      ATTR       �   �   &                  �   &  com.apple.quarantine q/0001;58880409;Microsoft\x20Outlook; 