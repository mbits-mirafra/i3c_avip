module mgc_ace_master_hdl #(
   int ADDR_WIDTH  = 64,
   int RDATA_WIDTH = 1024,
   int WDATA_WIDTH = 1024,
   int ID_WIDTH    = 30,
   int USER_WIDTH  = 4,
   int REGION_MAP_SIZE = 16,
   int SNOOP_DATA_WIDTH = 1024,
   int CACHE_LINE_SIZE = 7,
   string VIP_IF_UVM_NAME,
   string VIP_IF_UVM_CONTEXT,
   int snoop_data_channel_phase_BUFFER_MAX_ELEMENTS = 17, 
   int write_channel_phase_BUFFER_MAX_ELEMENTS = 17, 
   int BURST_BUFFER = 16,
   type PARAMS = int
)(mgc_ace_signal_if pin_if); //pragma attribute mgc_ace_master_hdl partition_module_xrtl

`ifdef XRTL

   //
   // Instantiate VTL XRTL BFM:
   //
   mgc_xrtl_ace_master #(
      .AXI4_ADDRESS_WIDTH(ADDR_WIDTH),
      .AXI4_RDATA_WIDTH(RDATA_WIDTH),
      .AXI4_WDATA_WIDTH(WDATA_WIDTH),
      .AXI4_ID_WIDTH(ID_WIDTH),
      .AXI4_USER_WIDTH(USER_WIDTH),
      .AXI4_REGION_MAP_SIZE(REGION_MAP_SIZE),
      .ACE_SNOOP_DATA_WIDTH(SNOOP_DATA_WIDTH),
      .ACE_CACHE_LINE_SIZE(CACHE_LINE_SIZE),
      .snoop_data_channel_phase_BUFFER_MAX_ELEMENTS(snoop_data_channel_phase_BUFFER_MAX_ELEMENTS),
      .write_channel_phase_BUFFER_MAX_ELEMENTS(write_channel_phase_BUFFER_MAX_ELEMENTS),
      .BURST_BUFFER(BURST_BUFFER)
   ) vip_module (
      .ACVALID(pin_if.ACVALID),
      .ACREADY(pin_if.ACREADY),
      .ACADDR(pin_if.ACADDR),
      .ACSNOOP(pin_if.ACSNOOP),
      .ACPROT(pin_if.ACPROT),
      .CDVALID(pin_if.CDVALID),
      .CDREADY(pin_if.CDREADY),
      .CDDATA(pin_if.CDDATA),
      .CDLAST(pin_if.CDLAST),
      .CRVALID(pin_if.CRVALID),
      .CRREADY(pin_if.CRREADY),
      .CRRESP(pin_if.CRRESP),
      .ACLK(pin_if.ACLK),
      .ARESETn(pin_if.ARESETn),
      .AWVALID(pin_if.AWVALID),
      .AWADDR(pin_if.AWADDR),
      .AWPROT(pin_if.AWPROT),
      .AWREGION(pin_if.AWREGION),
      .AWLEN(pin_if.AWLEN),
      .AWSIZE(pin_if.AWSIZE),
      .AWBURST(pin_if.AWBURST),
      .AWLOCK(pin_if.AWLOCK),
      .AWCACHE(pin_if.AWCACHE),
      .AWQOS(pin_if.AWQOS),
      .AWID(pin_if.AWID),
      .AWUSER(pin_if.AWUSER),
      .AWDOMAIN(pin_if.AWDOMAIN),
      .AWSNOOP(pin_if.AWSNOOP),
      .AWBAR(pin_if.AWBAR),
      .ARDOMAIN(pin_if.ARDOMAIN),
      .ARSNOOP(pin_if.ARSNOOP),
      .ARBAR(pin_if.ARBAR),
      .RRESP(pin_if.RRESP),
      .RACK(pin_if.RACK),
      .WACK(pin_if.WACK),
      .AWREADY(pin_if.AWREADY),
      .ARVALID(pin_if.ARVALID),
      .ARADDR(pin_if.ARADDR),
      .ARPROT(pin_if.ARPROT),
      .ARREGION(pin_if.ARREGION),
      .ARLEN(pin_if.ARLEN),
      .ARSIZE(pin_if.ARSIZE),
      .ARBURST(pin_if.ARBURST),
      .ARLOCK(pin_if.ARLOCK),
      .ARCACHE(pin_if.ARCACHE),
      .ARQOS(pin_if.ARQOS),
      .ARID(pin_if.ARID),
      .ARUSER(pin_if.ARUSER),
      .ARREADY(pin_if.ARREADY),
      .RVALID(pin_if.RVALID),
      .RDATA(pin_if.RDATA),
      .RLAST(pin_if.RLAST),
      .RID(pin_if.RID),
      .RUSER(pin_if.RUSER),
      .RREADY(pin_if.RREADY),
      .WVALID(pin_if.WVALID),
      .WDATA(pin_if.WDATA),
      .WSTRB(pin_if.WSTRB),
      .WLAST(pin_if.WLAST),
      .WUSER(pin_if.WUSER),
      .WREADY(pin_if.WREADY),
      .BVALID(pin_if.BVALID),
      .BRESP(pin_if.BRESP),
      .BID(pin_if.BID),
      .BUSER(pin_if.BUSER),
      .BREADY(pin_if.BREADY)
   );

`else

   //
   // Instantiate QVIP connectivity module:
   //
   ace_master #(
      .PARAMS(PARAMS),
      .IF_NAME(VIP_IF_UVM_NAME),
      .PATH_NAME(VIP_IF_UVM_CONTEXT)
   ) vip_module (
      .ACLK(pin_if.ACLK),
      .ARESETn(pin_if.ARESETn),
      .AWID(pin_if.AWID),
      .AWADDR(pin_if.AWADDR),
      .AWLEN(pin_if.AWLEN),
      .AWSIZE(pin_if.AWSIZE),
      .AWBURST(pin_if.AWBURST),
      .AWLOCK(pin_if.AWLOCK),
      .AWCACHE(pin_if.AWCACHE),
      .AWPROT(pin_if.AWPROT),
      .AWQOS(pin_if.AWQOS),
      .AWREGION(pin_if.AWREGION),
      .AWUSER(pin_if.AWUSER),
      .AWVALID(pin_if.AWVALID),
      .AWREADY(pin_if.AWREADY),
      .AWSNOOP(pin_if.AWSNOOP),
      .AWDOMAIN(pin_if.AWDOMAIN),
      .AWBAR(pin_if.AWBAR),
      .AWUNIQUE(pin_if.AWUNIQUE),
      .WDATA(pin_if.WDATA),
      .WSTRB(pin_if.WSTRB),
      .WLAST(pin_if.WLAST),
      .WUSER(pin_if.WUSER),
      .WVALID(pin_if.WVALID),
      .WREADY(pin_if.WREADY),
      .BID(pin_if.BID),
      .BRESP(pin_if.BRESP),
      .BUSER(pin_if.BUSER),
      .BVALID(pin_if.BVALID),
      .BREADY(pin_if.BREADY),
      .WACK(pin_if.WACK),
      .ARID(pin_if.ARID),
      .ARADDR(pin_if.ARADDR),
      .ARLEN(pin_if.ARLEN),
      .ARSIZE(pin_if.ARSIZE),
      .ARBURST(pin_if.ARBURST),
      .ARLOCK(pin_if.ARLOCK),
      .ARCACHE(pin_if.ARCACHE),
      .ARPROT(pin_if.ARPROT),
      .ARQOS(pin_if.ARQOS),
      .ARREGION(pin_if.ARREGION),
      .ARUSER(pin_if.ARUSER),
      .ARVALID(pin_if.ARVALID),
      .ARREADY(pin_if.ARREADY),
      .ARSNOOP(pin_if.ARSNOOP),
      .ARDOMAIN(pin_if.ARDOMAIN),
      .ARBAR(pin_if.ARBAR),
      .RID(pin_if.RID),
      .RDATA(pin_if.RDATA),
      .RRESP(pin_if.RRESP),
      .RLAST(pin_if.RLAST),
      .RUSER(pin_if.RUSER),
      .RVALID(pin_if.RVALID),
      .RREADY(pin_if.RREADY),
      .RACK(pin_if.RACK),
      .ACVALID(pin_if.ACVALID),
      .ACREADY(pin_if.ACREADY),
      .ACADDR(pin_if.ACADDR),
      .ACSNOOP(pin_if.ACSNOOP),
      .ACPROT(pin_if.ACPROT),
      .CRVALID(pin_if.CRVALID),
      .CRREADY(pin_if.CRREADY),
      .CRRESP(pin_if.CRRESP),
      .CDVALID(pin_if.CDVALID),
      .CDREADY(pin_if.CDREADY),
      .CDDATA(pin_if.CDDATA),
      .CDLAST(pin_if.CDLAST)
	 );

`endif

endmodule: mgc_ace_master_hdl
