//----------------------------------------------------------------------
// Created with uvmf_gen version 2019.4_1
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This file contains macros used with the alu_in package.
//   These macros include packed struct definitions.  These structs are
//   used to pass data between classes, hvl, and BFM's, hdl.  Use of 
//   structs are more efficient and simpler to modify.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_struct
//      and from_struct methods defined in the macros below that are used in  
//      the alu_in_configuration class.
//
  `define alu_in_CONFIGURATION_STRUCT \
typedef struct packed  { \
     uvmf_active_passive_t active_passive; \
     uvmf_initiator_responder_t initiator_responder; \
     } alu_in_configuration_s;

  `define alu_in_CONFIGURATION_TO_STRUCT_FUNCTION \
  virtual function alu_in_configuration_s to_struct();\
    alu_in_configuration_struct = \
       {\
       this.active_passive,\
       this.initiator_responder\
       };\
    return ( alu_in_configuration_struct );\
  endfunction

  `define alu_in_CONFIGURATION_FROM_STRUCT_FUNCTION \
  virtual function void from_struct(alu_in_configuration_s alu_in_configuration_struct);\
      {\
      this.active_passive,\
      this.initiator_responder  \
      } = alu_in_configuration_struct;\
  endfunction

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_monitor_struct
//      and from_monitor_struct methods of the alu_in_transaction class.
//
  `define alu_in_MONITOR_STRUCT typedef struct packed  { \
  alu_in_op_t op ; \
  bit [ALU_IN_OP_WIDTH-1:0] a ; \
  bit [ALU_IN_OP_WIDTH-1:0] b ; \
     } alu_in_monitor_s;

  `define alu_in_TO_MONITOR_STRUCT_FUNCTION \
  virtual function alu_in_monitor_s to_monitor_struct();\
    alu_in_monitor_struct = \
            { \
            this.op , \
            this.a , \
            this.b  \
            };\
    return ( alu_in_monitor_struct);\
  endfunction\

  `define alu_in_FROM_MONITOR_STRUCT_FUNCTION \
  virtual function void from_monitor_struct(alu_in_monitor_s alu_in_monitor_struct);\
            {\
            this.op , \
            this.a , \
            this.b  \
            } = alu_in_monitor_struct;\
  endfunction

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_initiator_struct
//      and from_initiator_struct methods of the alu_in_transaction class.
//      Also update the comments in the driver BFM.
//
  `define alu_in_INITIATOR_STRUCT typedef struct packed  { \
  alu_in_op_t op ; \
  bit [ALU_IN_OP_WIDTH-1:0] a ; \
  bit [ALU_IN_OP_WIDTH-1:0] b ; \
     } alu_in_initiator_s;

  `define alu_in_TO_INITIATOR_STRUCT_FUNCTION \
  virtual function alu_in_initiator_s to_initiator_struct();\
    alu_in_initiator_struct = \
           {\
           this.op , \
           this.a , \
           this.b  \
           };\
    return ( alu_in_initiator_struct);\
  endfunction

  `define alu_in_FROM_INITIATOR_STRUCT_FUNCTION \
  virtual function void from_initiator_struct(alu_in_initiator_s alu_in_initiator_struct);\
           {\
           this.op , \
           this.a , \
           this.b  \
           } = alu_in_initiator_struct;\
  endfunction

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_responder_struct
//      and from_responder_struct methods of the alu_in_transaction class.
//      Also update the comments in the driver BFM.
//
  `define alu_in_RESPONDER_STRUCT typedef struct packed  { \
  alu_in_op_t op ; \
  bit [ALU_IN_OP_WIDTH-1:0] a ; \
  bit [ALU_IN_OP_WIDTH-1:0] b ; \
     } alu_in_responder_s;

  `define alu_in_TO_RESPONDER_STRUCT_FUNCTION \
  virtual function alu_in_responder_s to_responder_struct();\
    alu_in_responder_struct = \
           {\
           this.op , \
           this.a , \
           this.b  \
           };\
    return ( alu_in_responder_struct);\
  endfunction

  `define alu_in_FROM_RESPONDER_STRUCT_FUNCTION \
  virtual function void from_responder_struct(alu_in_responder_s alu_in_responder_struct);\
           {\
           this.op , \
           this.a , \
           this.b  \
           } = alu_in_responder_struct;\
  endfunction
// pragma uvmf custom additional begin
// pragma uvmf custom additional end
