//
// File: test_packages.svh
//
// Generated from Mentor VIP Configurator (20200115)
// Generated using Mentor VIP Library ( 2020.1 : 01/23/2020:13:29 )
//

import qvip_agents_pkg::*;

// Add other packages here as required
