//
// File: test_packages.svh
//
// Generated from Mentor VIP Configurator (20160818)
// Generated using Mentor VIP Library ( 10_5b : 09/04/2016:09:24 )
//

import axi4_2x2_fabric_qvip_pkg::*;

// Add other packages here as required
