//
// File: qvip_agents_pkg.sv
//
// Generated from Mentor VIP Configurator (20200115)
// Generated using Mentor VIP Library ( 2020.1 : 01/23/2020:13:29 )
//
package qvip_agents_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    
    import addr_map_pkg::*;
    
    import qvip_agents_params_pkg::*;
    import mvc_pkg::*;
    import mgc_apb3_v1_0_pkg::*;
    
    `include "qvip_agents_env_config.svh"
    `include "qvip_agents_env.svh"
    `include "qvip_agents_vseq_base.svh"
    `include "qvip_agents_test_base.svh"
endpackage: qvip_agents_pkg
