//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// PACKAGE: This file defines all of the files contained in the
//    environment package that will run on the host simulator.
//
// CONTAINS:
//     - <env_configuration.svh>
//     - <env_environment.svh>
//     - <env_env_sequence_base.svh>
//     - <i3c_scoreboard.svh>
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
package env_env_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import uvmf_base_pkg::*;
  import i3c_m_pkg::*;
  import i3c_m_pkg_hdl::*;
  import i3c_s_pkg::*;
  import i3c_s_pkg_hdl::*;
 
  `uvm_analysis_imp_decl(_m_sb_ep)
  `uvm_analysis_imp_decl(_s_sb_ep)

  // pragma uvmf custom package_imports_additional begin
  // pragma uvmf custom package_imports_additional end

  // Parameters defined as HVL parameters

  `include "src/env_env_typedefs.svh"
  `include "src/env_env_configuration.svh"
  `include "src/i3c_scoreboard.svh"
  `include "src/env_environment.svh"
  `include "src/env_env_sequence_base.svh"

  // pragma uvmf custom package_item_additional begin
  // UVMF_CHANGE_ME : When adding new environment level sequences to the src directory
  //    be sure to add the sequence file here so that it will be
  //    compiled as part of the environment package.  Be sure to place
  //    the new sequence after any base sequence of the new sequence.
  // pragma uvmf custom package_item_additional end

endpackage

// pragma uvmf custom external begin
// pragma uvmf custom external end

