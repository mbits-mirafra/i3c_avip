//----------------------------------------------------------------------
// Created with uvmf_gen version 2020.1
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
// Description: This top level UVM test is the base class for all
//     future tests created for this project.
//
//     This test class contains:
//          Configuration:  The top level configuration for the project.
//          Environment:    The top level environment for the project.
//          Top_level_sequence:  The top level sequence for the project.
//                                        
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

typedef alu_env_configuration #(
        .APB_RDATA_WIDTH(TEST_APB_RDATA_WIDTH),
        .APB_WDATA_WIDTH(TEST_APB_WDATA_WIDTH),
        .APB_ADDR_WIDTH(TEST_APB_ADDR_WIDTH),
        .ALU_OUT_RESULT_WIDTH(TEST_ALU_OUT_RESULT_WIDTH),
        .ALU_IN_OP_WIDTH(TEST_ALU_IN_OP_WIDTH)
        )alu_env_configuration_t;
typedef alu_environment #(
        .APB_RDATA_WIDTH(TEST_APB_RDATA_WIDTH),
        .APB_WDATA_WIDTH(TEST_APB_WDATA_WIDTH),
        .APB_ADDR_WIDTH(TEST_APB_ADDR_WIDTH),
        .ALU_OUT_RESULT_WIDTH(TEST_ALU_OUT_RESULT_WIDTH),
        .ALU_IN_OP_WIDTH(TEST_ALU_IN_OP_WIDTH)
        )alu_environment_t;

class test_top extends uvmf_test_base #(.CONFIG_T(alu_env_configuration_t), 
                                        .ENV_T(alu_environment_t), 
                                        .TOP_LEVEL_SEQ_T(alu_bench_sequence_base));

  `uvm_component_utils( test_top );


  string interface_names[] = {
    uvm_test_top_environment_qvip_agents_env_apb_master_0 /* apb_master_0     [0] */ , 
    alu_in_agent_BFM /* alu_in_agent     [1] */ , 
    alu_out_agent_BFM /* alu_out_agent     [2] */ 
};

uvmf_active_passive_t interface_activities[] = { 
    ACTIVE /* apb_master_0     [0] */ , 
    ACTIVE /* alu_in_agent     [1] */ , 
    PASSIVE /* alu_out_agent     [2] */   };

  // pragma uvmf custom class_item_additional begin
  // pragma uvmf custom class_item_additional end

  // ****************************************************************************
  // FUNCTION: new()
  // This is the standard system verilog constructor.  All components are 
  // constructed in the build_phase to allow factory overriding.
  //
  function new( string name = "", uvm_component parent = null );
     super.new( name ,parent );
  endfunction



  // ****************************************************************************
  // FUNCTION: build_phase()
  // The construction of the configuration and environment classes is done in
  // the build_phase of uvmf_test_base.  Once the configuraton and environment
  // classes are built then the initialize call is made to perform the
  // following: 
  //     Monitor and driver BFM virtual interface handle passing into agents
  //     Set the active/passive state for each agent
  // Once this build_phase completes, the build_phase of the environment is
  // executed which builds the agents.
  //
  virtual function void build_phase(uvm_phase phase);

    // Turn on coverage for the Register Model
    uvm_reg::include_coverage("*", UVM_CVR_ALL);

    super.build_phase(phase);
    // pragma uvmf custom configuration_settings_post_randomize begin
    // pragma uvmf custom configuration_settings_post_randomize end
    configuration.initialize(NA, "uvm_test_top.environment", interface_names, null, interface_activities);
  endfunction

endclass
