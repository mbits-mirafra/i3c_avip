//----------------------------------------------------------------------
//   Copyright 2013 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------
//============================================================================
// @(#) $Id: XlSvTimeSync.svh 681 2011-07-06 10:56:19Z jstickle $
//============================================================================

`ifndef _XlSvTimeSync_svh_ // {
`define _XlSvTimeSync_svh_

//____________________                                       ________________
// class XlSvTimeSync \_____________________________________/ johnS 6-15-2010
//---------------------------------------------------------------------------

class XlSvTimeSync; // {

  //private:
    local event dIsAdvanceDone;
    local longint unsigned dScheduledClock;

  //public:

    function new(); endfunction

    //---------------------------------------------------------
    // accessors

    function void setScheduledClock( longint unsigned scheduledClock );
        dScheduledClock = scheduledClock; endfunction
    function longint unsigned scheduledClock();
        scheduledClock = dScheduledClock; endfunction

    task waitForSync(); @dIsAdvanceDone; endtask
    function void post(); ->dIsAdvanceDone; endfunction

  function string sprint();
    return $sformatf("dScheduledClock: %0d", dScheduledClock);
  endfunction : sprint
  
endclass // }

`endif // } _XlSvTimeSync_svh_
