//
// File: test_packages.svh
//
// Generated from Mentor VIP Configurator (20191003)
// Generated using Mentor VIP Library ( 2019.4 : 10/16/2019:13:47 )
//

import axi4_2x2_fabric_qvip_pkg::*;

// Add other packages here as required
