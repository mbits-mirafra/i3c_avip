//----------------------------------------------------------------------
// Created with uvmf_gen version 2021.1
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef enum bit[2:0] {CCS = 3'b000, CCS_RDY = 3'b001, CCS_VLD = 3'b010, CCS_WAIT = 3'b011, CCS_SYNC = 3'b100} protocol_kind_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

