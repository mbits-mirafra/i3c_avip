//
// File: axi4_2x2_fabric_qvip_pkg.sv
//
// Generated from Mentor VIP Configurator (20191003)
// Generated using Mentor VIP Library ( 2019.4 : 10/16/2019:13:47 )
//
package axi4_2x2_fabric_qvip_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    
    import addr_map_pkg::*;
    
    import axi4_2x2_fabric_qvip_params_pkg::*;
    import mvc_pkg::*;
    import mgc_axi4_v1_0_pkg::*;
    
    `include "axi4_2x2_fabric_qvip_env_config.svh"
    `include "axi4_2x2_fabric_qvip_env.svh"
    `include "axi4_2x2_fabric_qvip_vseq_base.svh"
    `include "axi4_2x2_fabric_qvip_test_base.svh"
endpackage: axi4_2x2_fabric_qvip_pkg
