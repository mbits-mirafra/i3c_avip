
//------> /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/pkgs/siflibs/ccs_conn_in_wait_v1.v 
module ccs_conn_in_wait_v1 (
  vld, rdy, dat, idat, irdy, ivld, clk, en, arst, srst
);

  parameter integer width = 32;
  parameter integer ph_clk  = 1;
  parameter integer ph_en   = 1;
  parameter integer ph_arst = 1;
  parameter integer ph_srst = 1;
  //parameter         has_en  = 1'b1;
  input [width-1:0] dat;
  input vld;
  output rdy;
  output [width-1:0] idat;
  input irdy;
  output ivld;
  input clk;
  input en;
  input arst;
  input srst;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld; 
endmodule




//------> /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/pkgs/siflibs/ccs_conn_out_wait_v1.v 
module ccs_conn_out_wait_v1 (
  vld, rdy, dat, idat, ivld, irdy,
      clk, en, arst, srst
);
  parameter integer width = 32;
  parameter integer ph_clk  = 1;
  parameter integer ph_en  = 1;
  parameter integer ph_arst = 1;
  parameter integer ph_srst = 1;
  //parameter         has_en  = 1'b1;
  output [width-1:0] dat;
  output vld;
  input rdy;
  input [width-1:0] idat;
  input ivld;
  output irdy;
  input clk;
  input en;
  input arst;
  input srst;
  
  assign dat = idat;
  assign vld = ivld;
  assign irdy = rdy; 

endmodule




//------> /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/pkgs/siflibs/ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ../td_ccore_solutions/Connections__Combinational_bool_Connections__SYN_PORT___Push_eb3219e1ee4a808220eaf5e336d914dd5e91_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6/912629 Production Release
//  HLS Date:       Thu Dec  3 18:37:23 PST 2020
// 
//  Generated by:   daerne@orw-lehavre-r77
//  Generated date: Wed Dec 16 18:35:46 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_bool_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_Combinational_bool_Connections_SYN_PORT_Push_core (
  this_vld, this_rdy, this_dat, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output this_dat;
  reg this_dat;
  input m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd1)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd89),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd97)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_3_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 1'b0;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_bool_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_Combinational_bool_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output this_dat;
  input m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_bool_Connections_SYN_PORT_Push_core Connections_Combinational_bool_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ../td_ccore_solutions/Connections__Combinational_bool_Connections__SYN_PORT___Pop_705d86a2cfe12487109e329e5525b57f5cfb_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6/912629 Production Release
//  HLS Date:       Thu Dec  3 18:37:23 PST 2020
// 
//  Generated by:   daerne@orw-lehavre-r77
//  Generated date: Wed Dec 16 18:35:44 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_bool_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module Connections_Combinational_bool_Connections_SYN_PORT_Pop_core (
  this_vld, this_rdy, this_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_2_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire  nl_return_rsci_d;
  assign nl_return_rsci_d = this_dat;
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_vld;
  mgc_out_dreg_v2 #(.rscid(32'sd12),
  .width(32'sd1)) return_rsci (
      .d(nl_return_rsci_d),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd88),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd96)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_2_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_vld));
  assign this_rdy_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_vld
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( or_2_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_2_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_bool_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module Connections_Combinational_bool_Connections_SYN_PORT_Pop (
  this_vld, this_rdy, this_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_bool_Connections_SYN_PORT_Pop_core Connections_Combinational_bool_Connections_SYN_PORT_Pop_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_dma_cmd_Connections__SYN_PORT__--_60d0a04a3fd75a59153aaacf532596ed899d_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6/912629 Production Release
//  HLS Date:       Thu Dec  3 18:37:23 PST 2020
// 
//  Generated by:   daerne@orw-lehavre-r77
//  Generated date: Tue Jan  5 16:52:07 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_dma_cmd_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_Combinational_dma_cmd_Connections_SYN_PORT_Push_core (
  this_vld, this_rdy, this_dat, m_ar_addr_rsc_dat, m_aw_addr_rsc_dat, m_total_len_rsc_dat,
      m_scatter_stride_rsc_dat, m_scatter_len_rsc_dat, m_scatter_groups_rsc_dat,
      m_dma_mode_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [175:0] this_dat;
  input [31:0] m_ar_addr_rsc_dat;
  input [31:0] m_aw_addr_rsc_dat;
  input [31:0] m_total_len_rsc_dat;
  input [31:0] m_scatter_stride_rsc_dat;
  input [15:0] m_scatter_len_rsc_dat;
  input [15:0] m_scatter_groups_rsc_dat;
  input [15:0] m_dma_mode_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [31:0] m_ar_addr_rsci_idat;
  wire [31:0] m_aw_addr_rsci_idat;
  wire [31:0] m_total_len_rsci_idat;
  wire [31:0] m_scatter_stride_rsci_idat;
  wire [15:0] m_scatter_len_rsci_idat;
  wire [15:0] m_scatter_groups_rsci_idat;
  wire [15:0] m_dma_mode_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [15:0] m_dma_mode_buf_lpi_1_dfm;
  reg [15:0] m_scatter_groups_buf_lpi_1_dfm;
  reg [15:0] m_scatter_len_buf_lpi_1_dfm;
  reg [31:0] m_scatter_stride_buf_lpi_1_dfm;
  reg [31:0] m_total_len_buf_lpi_1_dfm;
  reg [31:0] m_aw_addr_buf_lpi_1_dfm;
  reg [31:0] m_ar_addr_buf_lpi_1_dfm;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd38),
  .width(32'sd32)) m_ar_addr_rsci (
      .dat(m_ar_addr_rsc_dat),
      .idat(m_ar_addr_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd39),
  .width(32'sd32)) m_aw_addr_rsci (
      .dat(m_aw_addr_rsc_dat),
      .idat(m_aw_addr_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd40),
  .width(32'sd32)) m_total_len_rsci (
      .dat(m_total_len_rsc_dat),
      .idat(m_total_len_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd41),
  .width(32'sd32)) m_scatter_stride_rsci (
      .dat(m_scatter_stride_rsc_dat),
      .idat(m_scatter_stride_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd42),
  .width(32'sd16)) m_scatter_len_rsci (
      .dat(m_scatter_len_rsc_dat),
      .idat(m_scatter_len_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd43),
  .width(32'sd16)) m_scatter_groups_rsci (
      .dat(m_scatter_groups_rsc_dat),
      .idat(m_scatter_groups_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd44),
  .width(32'sd16)) m_dma_mode_rsci (
      .dat(m_dma_mode_rsc_dat),
      .idat(m_dma_mode_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd87),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd95)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = {m_dma_mode_buf_lpi_1_dfm , m_scatter_groups_buf_lpi_1_dfm ,
      m_scatter_len_buf_lpi_1_dfm , m_scatter_stride_buf_lpi_1_dfm , m_total_len_buf_lpi_1_dfm
      , m_aw_addr_buf_lpi_1_dfm , m_ar_addr_buf_lpi_1_dfm};
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_3_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_dma_mode_buf_lpi_1_dfm <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_dma_mode_buf_lpi_1_dfm <= m_dma_mode_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_scatter_groups_buf_lpi_1_dfm <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_scatter_groups_buf_lpi_1_dfm <= m_scatter_groups_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_scatter_len_buf_lpi_1_dfm <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_scatter_len_buf_lpi_1_dfm <= m_scatter_len_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_scatter_stride_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_scatter_stride_buf_lpi_1_dfm <= m_scatter_stride_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_total_len_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_total_len_buf_lpi_1_dfm <= m_total_len_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_aw_addr_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_aw_addr_buf_lpi_1_dfm <= m_aw_addr_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_ar_addr_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_ar_addr_buf_lpi_1_dfm <= m_ar_addr_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_dma_cmd_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_Combinational_dma_cmd_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_ar_addr_rsc_dat, m_aw_addr_rsc_dat, m_total_len_rsc_dat,
      m_scatter_stride_rsc_dat, m_scatter_len_rsc_dat, m_scatter_groups_rsc_dat,
      m_dma_mode_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [175:0] this_dat;
  input [31:0] m_ar_addr_rsc_dat;
  input [31:0] m_aw_addr_rsc_dat;
  input [31:0] m_total_len_rsc_dat;
  input [31:0] m_scatter_stride_rsc_dat;
  input [15:0] m_scatter_len_rsc_dat;
  input [15:0] m_scatter_groups_rsc_dat;
  input [15:0] m_dma_mode_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_dma_cmd_Connections_SYN_PORT_Push_core Connections_Combinational_dma_cmd_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_ar_addr_rsc_dat(m_ar_addr_rsc_dat),
      .m_aw_addr_rsc_dat(m_aw_addr_rsc_dat),
      .m_total_len_rsc_dat(m_total_len_rsc_dat),
      .m_scatter_stride_rsc_dat(m_scatter_stride_rsc_dat),
      .m_scatter_len_rsc_dat(m_scatter_len_rsc_dat),
      .m_scatter_groups_rsc_dat(m_scatter_groups_rsc_dat),
      .m_dma_mode_rsc_dat(m_dma_mode_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_dma_cmd_Connections__SYN_PORT__--_cbe0c26edc75a386df5c7a6460f51cc589ba_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6/912629 Production Release
//  HLS Date:       Thu Dec  3 18:37:23 PST 2020
// 
//  Generated by:   daerne@orw-lehavre-r77
//  Generated date: Wed Dec 16 18:35:39 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_dma_cmd_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module Connections_Combinational_dma_cmd_Connections_SYN_PORT_Pop_core (
  this_vld, this_rdy, this_dat, return_ar_addr_rsc_z, return_aw_addr_rsc_z, return_total_len_rsc_z,
      return_scatter_stride_rsc_z, return_scatter_len_rsc_z, return_scatter_groups_rsc_z,
      return_dma_mode_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [175:0] this_dat;
  output [31:0] return_ar_addr_rsc_z;
  output [31:0] return_aw_addr_rsc_z;
  output [31:0] return_total_len_rsc_z;
  output [31:0] return_scatter_stride_rsc_z;
  output [15:0] return_scatter_len_rsc_z;
  output [15:0] return_scatter_groups_rsc_z;
  output [15:0] return_dma_mode_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_2_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_return_ar_addr_rsci_d;
  assign nl_return_ar_addr_rsci_d = this_dat[31:0];
  wire [31:0] nl_return_aw_addr_rsci_d;
  assign nl_return_aw_addr_rsci_d = this_dat[63:32];
  wire [31:0] nl_return_total_len_rsci_d;
  assign nl_return_total_len_rsci_d = this_dat[95:64];
  wire [31:0] nl_return_scatter_stride_rsci_d;
  assign nl_return_scatter_stride_rsci_d = this_dat[127:96];
  wire [15:0] nl_return_scatter_len_rsci_d;
  assign nl_return_scatter_len_rsci_d = this_dat[143:128];
  wire [15:0] nl_return_scatter_groups_rsci_d;
  assign nl_return_scatter_groups_rsci_d = this_dat[159:144];
  wire [15:0] nl_return_dma_mode_rsci_d;
  assign nl_return_dma_mode_rsci_d = this_dat[175:160];
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_vld;
  mgc_out_dreg_v2 #(.rscid(32'sd46),
  .width(32'sd32)) return_ar_addr_rsci (
      .d(nl_return_ar_addr_rsci_d[31:0]),
      .z(return_ar_addr_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd47),
  .width(32'sd32)) return_aw_addr_rsci (
      .d(nl_return_aw_addr_rsci_d[31:0]),
      .z(return_aw_addr_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd48),
  .width(32'sd32)) return_total_len_rsci (
      .d(nl_return_total_len_rsci_d[31:0]),
      .z(return_total_len_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd49),
  .width(32'sd32)) return_scatter_stride_rsci (
      .d(nl_return_scatter_stride_rsci_d[31:0]),
      .z(return_scatter_stride_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd50),
  .width(32'sd16)) return_scatter_len_rsci (
      .d(nl_return_scatter_len_rsci_d[15:0]),
      .z(return_scatter_len_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd51),
  .width(32'sd16)) return_scatter_groups_rsci (
      .d(nl_return_scatter_groups_rsci_d[15:0]),
      .z(return_scatter_groups_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd52),
  .width(32'sd16)) return_dma_mode_rsci (
      .d(nl_return_dma_mode_rsci_d[15:0]),
      .z(return_dma_mode_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd86),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd94)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_2_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_vld));
  assign this_rdy_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_vld
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( or_2_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_2_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_dma_cmd_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module Connections_Combinational_dma_cmd_Connections_SYN_PORT_Pop (
  this_vld, this_rdy, this_dat, return_ar_addr_rsc_z, return_aw_addr_rsc_z, return_total_len_rsc_z,
      return_scatter_stride_rsc_z, return_scatter_len_rsc_z, return_scatter_groups_rsc_z,
      return_dma_mode_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [175:0] this_dat;
  output [31:0] return_ar_addr_rsc_z;
  output [31:0] return_aw_addr_rsc_z;
  output [31:0] return_total_len_rsc_z;
  output [31:0] return_scatter_stride_rsc_z;
  output [15:0] return_scatter_len_rsc_z;
  output [15:0] return_scatter_groups_rsc_z;
  output [15:0] return_dma_mode_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_dma_cmd_Connections_SYN_PORT_Pop_core Connections_Combinational_dma_cmd_Connections_SYN_PORT_Pop_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .return_ar_addr_rsc_z(return_ar_addr_rsc_z),
      .return_aw_addr_rsc_z(return_aw_addr_rsc_z),
      .return_total_len_rsc_z(return_total_len_rsc_z),
      .return_scatter_stride_rsc_z(return_scatter_stride_rsc_z),
      .return_scatter_len_rsc_z(return_scatter_len_rsc_z),
      .return_scatter_groups_rsc_z(return_scatter_groups_rsc_z),
      .return_dma_mode_rsc_z(return_dma_mode_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_axi__axi4_segment_axi__cfg__sta--_ca82636619f0fa57f3aa71c27146deef77ee_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6/912629 Production Release
//  HLS Date:       Thu Dec  3 18:37:23 PST 2020
// 
//  Generated by:   daerne@orw-lehavre-r77
//  Generated date: Wed Dec 16 18:35:37 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_ar_payload_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_ar_payload_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_addr_rsc_dat, m_ex_len_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [75:0] this_dat;
  input [31:0] m_addr_rsc_dat;
  input [31:0] m_ex_len_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [31:0] m_addr_rsci_idat;
  wire [31:0] m_ex_len_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [31:0] m_ex_len_buf_lpi_1_dfm;
  reg [31:0] m_addr_buf_lpi_1_dfm;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd54),
  .width(32'sd32)) m_addr_rsci (
      .dat(m_addr_rsc_dat),
      .idat(m_addr_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd56),
  .width(32'sd32)) m_ex_len_rsci (
      .dat(m_ex_len_rsc_dat),
      .idat(m_ex_len_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd85),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd93)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = {m_ex_len_buf_lpi_1_dfm , 8'b00000000 , m_addr_buf_lpi_1_dfm
      , 4'b0000};
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_3_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_ex_len_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_ex_len_buf_lpi_1_dfm <= m_ex_len_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_addr_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_addr_buf_lpi_1_dfm <= m_addr_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_ar_payload_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_ar_payload_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_addr_rsc_dat, m_ex_len_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [75:0] this_dat;
  input [31:0] m_addr_rsc_dat;
  input [31:0] m_ex_len_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_ar_payload_Connections_SYN_PORT_Push_core
      Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_ar_payload_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_addr_rsc_dat(m_addr_rsc_dat),
      .m_ex_len_rsc_dat(m_ex_len_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_axi__axi4_segment_axi__cfg__sta--_17b736e90ec0a175ee935b87a3343a9d77ee_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6/912629 Production Release
//  HLS Date:       Thu Dec  3 18:37:23 PST 2020
// 
//  Generated by:   daerne@orw-lehavre-r77
//  Generated date: Wed Dec 16 18:35:35 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_aw_payload_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_aw_payload_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_addr_rsc_dat, m_ex_len_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [75:0] this_dat;
  input [31:0] m_addr_rsc_dat;
  input [31:0] m_ex_len_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [31:0] m_addr_rsci_idat;
  wire [31:0] m_ex_len_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [31:0] m_ex_len_buf_lpi_1_dfm;
  reg [31:0] m_addr_buf_lpi_1_dfm;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd58),
  .width(32'sd32)) m_addr_rsci (
      .dat(m_addr_rsc_dat),
      .idat(m_addr_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd60),
  .width(32'sd32)) m_ex_len_rsci (
      .dat(m_ex_len_rsc_dat),
      .idat(m_ex_len_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd84),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd92)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = {m_ex_len_buf_lpi_1_dfm , 8'b00000000 , m_addr_buf_lpi_1_dfm
      , 4'b0000};
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_3_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_ex_len_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_ex_len_buf_lpi_1_dfm <= m_ex_len_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_addr_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_addr_buf_lpi_1_dfm <= m_addr_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_aw_payload_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_aw_payload_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_addr_rsc_dat, m_ex_len_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [75:0] this_dat;
  input [31:0] m_addr_rsc_dat;
  input [31:0] m_ex_len_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_aw_payload_Connections_SYN_PORT_Push_core
      Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_aw_payload_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_addr_rsc_dat(m_addr_rsc_dat),
      .m_ex_len_rsc_dat(m_ex_len_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_axi__axi4_axi__cfg__standard___--_2df71452371de2d3d625bc078dfe011d6e5d_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6/912629 Production Release
//  HLS Date:       Thu Dec  3 18:37:23 PST 2020
// 
//  Generated by:   daerne@orw-lehavre-r77
//  Generated date: Wed Dec 16 18:35:33 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_Combinational_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [72:0] this_dat;
  input [63:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [63:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [63:0] m_data_buf_lpi_1_dfm;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  reg reg_510_1_reg_1;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd65),
  .width(32'sd64)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd83),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd91)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = signext_73_66({reg_510_1_reg_1 , 1'b0 , m_data_buf_lpi_1_dfm});
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      reg_510_1_reg_1 <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      reg_510_1_reg_1 <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_lpi_1_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      m_data_buf_lpi_1_dfm <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end

  function automatic [72:0] signext_73_66;
    input [65:0] vector;
  begin
    signext_73_66= {{7{vector[65]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_Combinational_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [72:0] this_dat;
  input [63:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_Push_core
      Connections_Combinational_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_axi__axi4_axi__cfg__standard___--_f19ea0f98d4a076d2a63665693c758bf6969_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6/912629 Production Release
//  HLS Date:       Thu Dec  3 18:37:23 PST 2020
// 
//  Generated by:   daerne@orw-lehavre-r77
//  Generated date: Wed Dec 16 18:35:31 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_axi_axi4_axi_cfg_standard_WRespPayload_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module Connections_Combinational_axi_axi4_axi_cfg_standard_WRespPayload_Connections_SYN_PORT_Pop_core
    (
  this_vld, this_rdy, this_dat, return_id_rsc_z, return_resp_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [5:0] this_dat;
  output [3:0] return_id_rsc_z;
  output [1:0] return_resp_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_2_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire [3:0] nl_return_id_rsci_d;
  assign nl_return_id_rsci_d = this_dat[3:0];
  wire [1:0] nl_return_resp_rsci_d;
  assign nl_return_resp_rsci_d = this_dat[5:4];
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_vld;
  mgc_out_dreg_v2 #(.rscid(32'sd68),
  .width(32'sd4)) return_id_rsci (
      .d(nl_return_id_rsci_d[3:0]),
      .z(return_id_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd69),
  .width(32'sd2)) return_resp_rsci (
      .d(nl_return_resp_rsci_d[1:0]),
      .z(return_resp_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd82),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd90)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_2_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_vld));
  assign this_rdy_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_vld
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( or_2_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_2_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_axi_axi4_axi_cfg_standard_WRespPayload_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module Connections_Combinational_axi_axi4_axi_cfg_standard_WRespPayload_Connections_SYN_PORT_Pop
    (
  this_vld, this_rdy, this_dat, return_id_rsc_z, return_resp_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [5:0] this_dat;
  output [3:0] return_id_rsc_z;
  output [1:0] return_resp_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_axi_axi4_axi_cfg_standard_WRespPayload_Connections_SYN_PORT_Pop_core
      Connections_Combinational_axi_axi4_axi_cfg_standard_WRespPayload_Connections_SYN_PORT_Pop_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .return_id_rsc_z(return_id_rsc_z),
      .return_resp_rsc_z(return_resp_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.6/912629 Production Release
//  HLS Date:       Thu Dec  3 18:37:23 PST 2020
// 
//  Generated by:   daerne@orw-lehavre-r77
//  Generated date: Thu Jan  7 15:08:39 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_master_process_fsm
//  FSM Module
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_master_process_fsm (
  clk, rst_bar, master_process_wen, fsm_output, while_C_2_tr0, while_C_2_tr1, while_C_2_tr2,
      while_case_0_while_C_0_tr0, while_case_1_while_while_C_0_tr0, while_case_1_while_C_3_tr0,
      while_case_2_while_while_C_0_tr0, while_case_2_while_C_2_tr0
);
  input clk;
  input rst_bar;
  input master_process_wen;
  output [16:0] fsm_output;
  reg [16:0] fsm_output;
  input while_C_2_tr0;
  input while_C_2_tr1;
  input while_C_2_tr2;
  input while_case_0_while_C_0_tr0;
  input while_case_1_while_while_C_0_tr0;
  input while_case_1_while_C_3_tr0;
  input while_case_2_while_while_C_0_tr0;
  input while_case_2_while_C_2_tr0;


  // FSM State Type Declaration for scatter_gather_dma_master_process_master_process_fsm_1
  parameter
    master_process_rlp_C_0 = 5'd0,
    while_C_0 = 5'd1,
    while_C_1 = 5'd2,
    while_C_2 = 5'd3,
    while_case_0_while_C_0 = 5'd4,
    while_case_1_while_C_0 = 5'd5,
    while_case_1_while_C_1 = 5'd6,
    while_case_1_while_while_C_0 = 5'd7,
    while_case_1_while_C_2 = 5'd8,
    while_case_1_while_C_3 = 5'd9,
    while_case_2_while_C_0 = 5'd10,
    while_case_2_while_C_1 = 5'd11,
    while_case_2_while_while_C_0 = 5'd12,
    while_case_2_while_C_2 = 5'd13,
    while_C_3 = 5'd14,
    while_C_4 = 5'd15,
    while_C_5 = 5'd16;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : scatter_gather_dma_master_process_master_process_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 17'b00000000000000010;
        state_var_NS = while_C_1;
      end
      while_C_1 : begin
        fsm_output = 17'b00000000000000100;
        state_var_NS = while_C_2;
      end
      while_C_2 : begin
        fsm_output = 17'b00000000000001000;
        if ( while_C_2_tr0 ) begin
          state_var_NS = while_C_3;
        end
        else if ( while_C_2_tr1 ) begin
          state_var_NS = while_case_0_while_C_0;
        end
        else if ( while_C_2_tr2 ) begin
          state_var_NS = while_case_1_while_C_0;
        end
        else begin
          state_var_NS = while_case_2_while_C_0;
        end
      end
      while_case_0_while_C_0 : begin
        fsm_output = 17'b00000000000010000;
        if ( while_case_0_while_C_0_tr0 ) begin
          state_var_NS = while_C_3;
        end
        else begin
          state_var_NS = while_case_0_while_C_0;
        end
      end
      while_case_1_while_C_0 : begin
        fsm_output = 17'b00000000000100000;
        state_var_NS = while_case_1_while_C_1;
      end
      while_case_1_while_C_1 : begin
        fsm_output = 17'b00000000001000000;
        state_var_NS = while_case_1_while_while_C_0;
      end
      while_case_1_while_while_C_0 : begin
        fsm_output = 17'b00000000010000000;
        if ( while_case_1_while_while_C_0_tr0 ) begin
          state_var_NS = while_case_1_while_C_2;
        end
        else begin
          state_var_NS = while_case_1_while_while_C_0;
        end
      end
      while_case_1_while_C_2 : begin
        fsm_output = 17'b00000000100000000;
        state_var_NS = while_case_1_while_C_3;
      end
      while_case_1_while_C_3 : begin
        fsm_output = 17'b00000001000000000;
        if ( while_case_1_while_C_3_tr0 ) begin
          state_var_NS = while_C_3;
        end
        else begin
          state_var_NS = while_case_1_while_C_0;
        end
      end
      while_case_2_while_C_0 : begin
        fsm_output = 17'b00000010000000000;
        state_var_NS = while_case_2_while_C_1;
      end
      while_case_2_while_C_1 : begin
        fsm_output = 17'b00000100000000000;
        state_var_NS = while_case_2_while_while_C_0;
      end
      while_case_2_while_while_C_0 : begin
        fsm_output = 17'b00001000000000000;
        if ( while_case_2_while_while_C_0_tr0 ) begin
          state_var_NS = while_case_2_while_C_2;
        end
        else begin
          state_var_NS = while_case_2_while_while_C_0;
        end
      end
      while_case_2_while_C_2 : begin
        fsm_output = 17'b00010000000000000;
        if ( while_case_2_while_C_2_tr0 ) begin
          state_var_NS = while_C_3;
        end
        else begin
          state_var_NS = while_case_2_while_C_0;
        end
      end
      while_C_3 : begin
        fsm_output = 17'b00100000000000000;
        state_var_NS = while_C_4;
      end
      while_C_4 : begin
        fsm_output = 17'b01000000000000000;
        state_var_NS = while_C_5;
      end
      while_C_5 : begin
        fsm_output = 17'b10000000000000000;
        state_var_NS = while_C_0;
      end
      // master_process_rlp_C_0
      default : begin
        fsm_output = 17'b00000000000000001;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      state_var <= master_process_rlp_C_0;
    end
    else if ( master_process_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_staller_1
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_staller_1 (
  clk, rst_bar, master_process_flen_unreg, master_process_wen, master_process_wten,
      dma_cmd_chan_Pop_mioi_wen_comp, r_segment0_ex_ar_chan_Push_mioi_wen_comp, w_segment0_ex_aw_chan_Push_mioi_wen_comp,
      r_master0_r_Pop_mioi_wen_comp, w_segment0_w_chan_Push_mioi_wen_comp, w_segment0_b_chan_Pop_mioi_wen_comp,
      dma_done_Push_mioi_wen_comp
);
  input clk;
  input rst_bar;
  input master_process_flen_unreg;
  output master_process_wen;
  output master_process_wten;
  input dma_cmd_chan_Pop_mioi_wen_comp;
  input r_segment0_ex_ar_chan_Push_mioi_wen_comp;
  input w_segment0_ex_aw_chan_Push_mioi_wen_comp;
  input r_master0_r_Pop_mioi_wen_comp;
  input w_segment0_w_chan_Push_mioi_wen_comp;
  input w_segment0_b_chan_Pop_mioi_wen_comp;
  input dma_done_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg master_process_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign master_process_wen = dma_cmd_chan_Pop_mioi_wen_comp & r_segment0_ex_ar_chan_Push_mioi_wen_comp
      & w_segment0_ex_aw_chan_Push_mioi_wen_comp & r_master0_r_Pop_mioi_wen_comp
      & w_segment0_w_chan_Push_mioi_wen_comp & w_segment0_b_chan_Pop_mioi_wen_comp
      & dma_done_Push_mioi_wen_comp & (~ master_process_flen_unreg);
  assign master_process_wten = master_process_wten_reg;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      master_process_wten_reg <= 1'b0;
    end
    else begin
      master_process_wten_reg <= ~ master_process_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_dma_done_Push_mioi_dma_done_Push_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_dma_done_Push_mioi_dma_done_Push_mio_wait_dp
    (
  clk, rst_bar, dma_done_Push_mioi_oswt, dma_done_Push_mioi_wen_comp, dma_done_Push_mioi_biwt,
      dma_done_Push_mioi_bdwt, dma_done_Push_mioi_bcwt
);
  input clk;
  input rst_bar;
  input dma_done_Push_mioi_oswt;
  output dma_done_Push_mioi_wen_comp;
  input dma_done_Push_mioi_biwt;
  input dma_done_Push_mioi_bdwt;
  output dma_done_Push_mioi_bcwt;
  reg dma_done_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_done_Push_mioi_wen_comp = (~ dma_done_Push_mioi_oswt) | dma_done_Push_mioi_biwt
      | dma_done_Push_mioi_bcwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      dma_done_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_done_Push_mioi_bcwt <= ~((~(dma_done_Push_mioi_bcwt | dma_done_Push_mioi_biwt))
          | dma_done_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_dma_done_Push_mioi_dma_done_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_dma_done_Push_mioi_dma_done_Push_mio_wait_ctrl
    (
  master_process_wen, dma_done_Push_mioi_oswt, dma_done_Push_mioi_biwt, dma_done_Push_mioi_bdwt,
      dma_done_Push_mioi_bcwt, dma_done_Push_mioi_idat_master_process_sct, dma_done_Push_mioi_irdy
);
  input master_process_wen;
  input dma_done_Push_mioi_oswt;
  output dma_done_Push_mioi_biwt;
  output dma_done_Push_mioi_bdwt;
  input dma_done_Push_mioi_bcwt;
  output dma_done_Push_mioi_idat_master_process_sct;
  input dma_done_Push_mioi_irdy;


  // Interconnect Declarations
  wire dma_done_Push_mioi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_done_Push_mioi_bdwt = dma_done_Push_mioi_oswt & master_process_wen;
  assign dma_done_Push_mioi_biwt = dma_done_Push_mioi_ogwt & dma_done_Push_mioi_irdy;
  assign dma_done_Push_mioi_ogwt = dma_done_Push_mioi_oswt & (~ dma_done_Push_mioi_bcwt);
  assign dma_done_Push_mioi_idat_master_process_sct = dma_done_Push_mioi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi_w_segment0_b_chan_Pop_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi_w_segment0_b_chan_Pop_mio_wait_dp
    (
  clk, rst_bar, w_segment0_b_chan_Pop_mioi_oswt, w_segment0_b_chan_Pop_mioi_wen_comp,
      w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt, w_segment0_b_chan_Pop_mioi_biwt,
      w_segment0_b_chan_Pop_mioi_bdwt, w_segment0_b_chan_Pop_mioi_bcwt, w_segment0_b_chan_Pop_mioi_return_resp_rsc_z
);
  input clk;
  input rst_bar;
  input w_segment0_b_chan_Pop_mioi_oswt;
  output w_segment0_b_chan_Pop_mioi_wen_comp;
  output [1:0] w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt;
  input w_segment0_b_chan_Pop_mioi_biwt;
  input w_segment0_b_chan_Pop_mioi_bdwt;
  output w_segment0_b_chan_Pop_mioi_bcwt;
  reg w_segment0_b_chan_Pop_mioi_bcwt;
  input [1:0] w_segment0_b_chan_Pop_mioi_return_resp_rsc_z;


  // Interconnect Declarations
  reg [1:0] w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_segment0_b_chan_Pop_mioi_wen_comp = (~ w_segment0_b_chan_Pop_mioi_oswt)
      | w_segment0_b_chan_Pop_mioi_biwt | w_segment0_b_chan_Pop_mioi_bcwt;
  assign w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt = MUX_v_2_2_2(w_segment0_b_chan_Pop_mioi_return_resp_rsc_z,
      w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_bfwt, w_segment0_b_chan_Pop_mioi_bcwt);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_segment0_b_chan_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      w_segment0_b_chan_Pop_mioi_bcwt <= ~((~(w_segment0_b_chan_Pop_mioi_bcwt | w_segment0_b_chan_Pop_mioi_biwt))
          | w_segment0_b_chan_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_bfwt <= 2'b00;
    end
    else if ( w_segment0_b_chan_Pop_mioi_biwt ) begin
      w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_bfwt <= w_segment0_b_chan_Pop_mioi_return_resp_rsc_z;
    end
  end

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi_w_segment0_b_chan_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi_w_segment0_b_chan_Pop_mio_wait_ctrl
    (
  master_process_wen, w_segment0_b_chan_Pop_mioi_oswt, w_segment0_b_chan_Pop_mioi_biwt,
      w_segment0_b_chan_Pop_mioi_bdwt, w_segment0_b_chan_Pop_mioi_bcwt, w_segment0_b_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct,
      w_segment0_b_chan_Pop_mioi_ccs_ccore_done_sync_vld, w_segment0_b_chan_Pop_mioi_oswt_pff
);
  input master_process_wen;
  input w_segment0_b_chan_Pop_mioi_oswt;
  output w_segment0_b_chan_Pop_mioi_biwt;
  output w_segment0_b_chan_Pop_mioi_bdwt;
  input w_segment0_b_chan_Pop_mioi_bcwt;
  output w_segment0_b_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  input w_segment0_b_chan_Pop_mioi_ccs_ccore_done_sync_vld;
  input w_segment0_b_chan_Pop_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign w_segment0_b_chan_Pop_mioi_bdwt = w_segment0_b_chan_Pop_mioi_oswt & master_process_wen;
  assign w_segment0_b_chan_Pop_mioi_biwt = w_segment0_b_chan_Pop_mioi_oswt & (~ w_segment0_b_chan_Pop_mioi_bcwt)
      & w_segment0_b_chan_Pop_mioi_ccs_ccore_done_sync_vld;
  assign w_segment0_b_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct =
      master_process_wen & w_segment0_b_chan_Pop_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_w_segment0_w_chan_Push_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_w_segment0_w_chan_Push_mio_wait_dp
    (
  clk, rst_bar, w_segment0_w_chan_Push_mioi_oswt_unreg, w_segment0_w_chan_Push_mioi_bawt,
      w_segment0_w_chan_Push_mioi_wen_comp, w_segment0_w_chan_Push_mioi_biwt, w_segment0_w_chan_Push_mioi_bdwt
);
  input clk;
  input rst_bar;
  input w_segment0_w_chan_Push_mioi_oswt_unreg;
  output w_segment0_w_chan_Push_mioi_bawt;
  output w_segment0_w_chan_Push_mioi_wen_comp;
  input w_segment0_w_chan_Push_mioi_biwt;
  input w_segment0_w_chan_Push_mioi_bdwt;


  // Interconnect Declarations
  reg w_segment0_w_chan_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_segment0_w_chan_Push_mioi_bawt = w_segment0_w_chan_Push_mioi_biwt | w_segment0_w_chan_Push_mioi_bcwt;
  assign w_segment0_w_chan_Push_mioi_wen_comp = (~ w_segment0_w_chan_Push_mioi_oswt_unreg)
      | w_segment0_w_chan_Push_mioi_bawt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_segment0_w_chan_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      w_segment0_w_chan_Push_mioi_bcwt <= ~((~(w_segment0_w_chan_Push_mioi_bcwt |
          w_segment0_w_chan_Push_mioi_biwt)) | w_segment0_w_chan_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_w_segment0_w_chan_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_w_segment0_w_chan_Push_mio_wait_ctrl
    (
  clk, rst_bar, w_segment0_w_chan_Push_mioi_oswt_unreg, master_process_wen, master_process_wten,
      w_segment0_w_chan_Push_mioi_iswt0, w_segment0_w_chan_Push_mioi_biwt, w_segment0_w_chan_Push_mioi_bdwt,
      w_segment0_w_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct, w_segment0_w_chan_Push_mioi_ccs_ccore_done_sync_vld,
      w_segment0_w_chan_Push_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  input w_segment0_w_chan_Push_mioi_oswt_unreg;
  input master_process_wen;
  input master_process_wten;
  input w_segment0_w_chan_Push_mioi_iswt0;
  output w_segment0_w_chan_Push_mioi_biwt;
  output w_segment0_w_chan_Push_mioi_bdwt;
  output w_segment0_w_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  input w_segment0_w_chan_Push_mioi_ccs_ccore_done_sync_vld;
  input w_segment0_w_chan_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire w_segment0_w_chan_Push_mioi_ogwt;
  reg w_segment0_w_chan_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_segment0_w_chan_Push_mioi_bdwt = w_segment0_w_chan_Push_mioi_oswt_unreg
      & master_process_wen;
  assign w_segment0_w_chan_Push_mioi_biwt = w_segment0_w_chan_Push_mioi_ogwt & w_segment0_w_chan_Push_mioi_ccs_ccore_done_sync_vld;
  assign w_segment0_w_chan_Push_mioi_ogwt = ((~ master_process_wten) & w_segment0_w_chan_Push_mioi_iswt0)
      | w_segment0_w_chan_Push_mioi_icwt;
  assign w_segment0_w_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct =
      master_process_wen & w_segment0_w_chan_Push_mioi_iswt0_pff;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_segment0_w_chan_Push_mioi_icwt <= 1'b0;
    end
    else begin
      w_segment0_w_chan_Push_mioi_icwt <= w_segment0_w_chan_Push_mioi_ogwt & (~ w_segment0_w_chan_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_r_master0_r_Pop_mioi_r_master0_r_Pop_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_r_master0_r_Pop_mioi_r_master0_r_Pop_mio_wait_dp
    (
  clk, rst_bar, r_master0_r_Pop_mioi_oswt_unreg, r_master0_r_Pop_mioi_bawt, r_master0_r_Pop_mioi_wen_comp,
      r_master0_r_Pop_mioi_idat_mxwt, r_master0_r_Pop_mioi_biwt, r_master0_r_Pop_mioi_bdwt,
      r_master0_r_Pop_mioi_idat
);
  input clk;
  input rst_bar;
  input r_master0_r_Pop_mioi_oswt_unreg;
  output r_master0_r_Pop_mioi_bawt;
  output r_master0_r_Pop_mioi_wen_comp;
  output [63:0] r_master0_r_Pop_mioi_idat_mxwt;
  input r_master0_r_Pop_mioi_biwt;
  input r_master0_r_Pop_mioi_bdwt;
  input [70:0] r_master0_r_Pop_mioi_idat;


  // Interconnect Declarations
  reg r_master0_r_Pop_mioi_bcwt;
  reg [63:0] r_master0_r_Pop_mioi_idat_bfwt_67_4;


  // Interconnect Declarations for Component Instantiations 
  assign r_master0_r_Pop_mioi_bawt = r_master0_r_Pop_mioi_biwt | r_master0_r_Pop_mioi_bcwt;
  assign r_master0_r_Pop_mioi_wen_comp = (~ r_master0_r_Pop_mioi_oswt_unreg) | r_master0_r_Pop_mioi_bawt;
  assign r_master0_r_Pop_mioi_idat_mxwt = MUX_v_64_2_2((r_master0_r_Pop_mioi_idat[67:4]),
      r_master0_r_Pop_mioi_idat_bfwt_67_4, r_master0_r_Pop_mioi_bcwt);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      r_master0_r_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      r_master0_r_Pop_mioi_bcwt <= ~((~(r_master0_r_Pop_mioi_bcwt | r_master0_r_Pop_mioi_biwt))
          | r_master0_r_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      r_master0_r_Pop_mioi_idat_bfwt_67_4 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( r_master0_r_Pop_mioi_biwt ) begin
      r_master0_r_Pop_mioi_idat_bfwt_67_4 <= r_master0_r_Pop_mioi_idat[67:4];
    end
  end

  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_r_master0_r_Pop_mioi_r_master0_r_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_r_master0_r_Pop_mioi_r_master0_r_Pop_mio_wait_ctrl
    (
  clk, rst_bar, r_master0_r_Pop_mioi_oswt_unreg, master_process_wen, master_process_wten,
      r_master0_r_Pop_mioi_iswt0, r_master0_r_Pop_mioi_biwt, r_master0_r_Pop_mioi_bdwt,
      r_master0_r_Pop_mioi_irdy_master_process_sct, r_master0_r_Pop_mioi_ivld
);
  input clk;
  input rst_bar;
  input r_master0_r_Pop_mioi_oswt_unreg;
  input master_process_wen;
  input master_process_wten;
  input r_master0_r_Pop_mioi_iswt0;
  output r_master0_r_Pop_mioi_biwt;
  output r_master0_r_Pop_mioi_bdwt;
  output r_master0_r_Pop_mioi_irdy_master_process_sct;
  input r_master0_r_Pop_mioi_ivld;


  // Interconnect Declarations
  wire r_master0_r_Pop_mioi_ogwt;
  reg r_master0_r_Pop_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign r_master0_r_Pop_mioi_bdwt = r_master0_r_Pop_mioi_oswt_unreg & master_process_wen;
  assign r_master0_r_Pop_mioi_biwt = r_master0_r_Pop_mioi_ogwt & r_master0_r_Pop_mioi_ivld;
  assign r_master0_r_Pop_mioi_ogwt = ((~ master_process_wten) & r_master0_r_Pop_mioi_iswt0)
      | r_master0_r_Pop_mioi_icwt;
  assign r_master0_r_Pop_mioi_irdy_master_process_sct = r_master0_r_Pop_mioi_ogwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      r_master0_r_Pop_mioi_icwt <= 1'b0;
    end
    else begin
      r_master0_r_Pop_mioi_icwt <= r_master0_r_Pop_mioi_ogwt & (~ r_master0_r_Pop_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_w_segment0_ex_aw_chan_Push_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_w_segment0_ex_aw_chan_Push_mio_wait_dp
    (
  clk, rst_bar, w_segment0_ex_aw_chan_Push_mioi_oswt, w_segment0_ex_aw_chan_Push_mioi_wen_comp,
      w_segment0_ex_aw_chan_Push_mioi_biwt, w_segment0_ex_aw_chan_Push_mioi_bdwt,
      w_segment0_ex_aw_chan_Push_mioi_bcwt
);
  input clk;
  input rst_bar;
  input w_segment0_ex_aw_chan_Push_mioi_oswt;
  output w_segment0_ex_aw_chan_Push_mioi_wen_comp;
  input w_segment0_ex_aw_chan_Push_mioi_biwt;
  input w_segment0_ex_aw_chan_Push_mioi_bdwt;
  output w_segment0_ex_aw_chan_Push_mioi_bcwt;
  reg w_segment0_ex_aw_chan_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign w_segment0_ex_aw_chan_Push_mioi_wen_comp = (~ w_segment0_ex_aw_chan_Push_mioi_oswt)
      | w_segment0_ex_aw_chan_Push_mioi_biwt | w_segment0_ex_aw_chan_Push_mioi_bcwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_segment0_ex_aw_chan_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      w_segment0_ex_aw_chan_Push_mioi_bcwt <= ~((~(w_segment0_ex_aw_chan_Push_mioi_bcwt
          | w_segment0_ex_aw_chan_Push_mioi_biwt)) | w_segment0_ex_aw_chan_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_w_segment0_ex_aw_chan_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_w_segment0_ex_aw_chan_Push_mio_wait_ctrl
    (
  master_process_wen, w_segment0_ex_aw_chan_Push_mioi_oswt, w_segment0_ex_aw_chan_Push_mioi_biwt,
      w_segment0_ex_aw_chan_Push_mioi_bdwt, w_segment0_ex_aw_chan_Push_mioi_bcwt,
      w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct,
      w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_done_sync_vld, w_segment0_ex_aw_chan_Push_mioi_oswt_pff
);
  input master_process_wen;
  input w_segment0_ex_aw_chan_Push_mioi_oswt;
  output w_segment0_ex_aw_chan_Push_mioi_biwt;
  output w_segment0_ex_aw_chan_Push_mioi_bdwt;
  input w_segment0_ex_aw_chan_Push_mioi_bcwt;
  output w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  input w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_done_sync_vld;
  input w_segment0_ex_aw_chan_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign w_segment0_ex_aw_chan_Push_mioi_bdwt = w_segment0_ex_aw_chan_Push_mioi_oswt
      & master_process_wen;
  assign w_segment0_ex_aw_chan_Push_mioi_biwt = w_segment0_ex_aw_chan_Push_mioi_oswt
      & (~ w_segment0_ex_aw_chan_Push_mioi_bcwt) & w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_done_sync_vld;
  assign w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct
      = master_process_wen & w_segment0_ex_aw_chan_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_r_segment0_ex_ar_chan_Push_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_r_segment0_ex_ar_chan_Push_mio_wait_dp
    (
  clk, rst_bar, r_segment0_ex_ar_chan_Push_mioi_oswt, r_segment0_ex_ar_chan_Push_mioi_wen_comp,
      r_segment0_ex_ar_chan_Push_mioi_biwt, r_segment0_ex_ar_chan_Push_mioi_bdwt,
      r_segment0_ex_ar_chan_Push_mioi_bcwt
);
  input clk;
  input rst_bar;
  input r_segment0_ex_ar_chan_Push_mioi_oswt;
  output r_segment0_ex_ar_chan_Push_mioi_wen_comp;
  input r_segment0_ex_ar_chan_Push_mioi_biwt;
  input r_segment0_ex_ar_chan_Push_mioi_bdwt;
  output r_segment0_ex_ar_chan_Push_mioi_bcwt;
  reg r_segment0_ex_ar_chan_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign r_segment0_ex_ar_chan_Push_mioi_wen_comp = (~ r_segment0_ex_ar_chan_Push_mioi_oswt)
      | r_segment0_ex_ar_chan_Push_mioi_biwt | r_segment0_ex_ar_chan_Push_mioi_bcwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      r_segment0_ex_ar_chan_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      r_segment0_ex_ar_chan_Push_mioi_bcwt <= ~((~(r_segment0_ex_ar_chan_Push_mioi_bcwt
          | r_segment0_ex_ar_chan_Push_mioi_biwt)) | r_segment0_ex_ar_chan_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_r_segment0_ex_ar_chan_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_r_segment0_ex_ar_chan_Push_mio_wait_ctrl
    (
  master_process_wen, r_segment0_ex_ar_chan_Push_mioi_oswt, r_segment0_ex_ar_chan_Push_mioi_biwt,
      r_segment0_ex_ar_chan_Push_mioi_bdwt, r_segment0_ex_ar_chan_Push_mioi_bcwt,
      r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct,
      r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_done_sync_vld, r_segment0_ex_ar_chan_Push_mioi_oswt_pff
);
  input master_process_wen;
  input r_segment0_ex_ar_chan_Push_mioi_oswt;
  output r_segment0_ex_ar_chan_Push_mioi_biwt;
  output r_segment0_ex_ar_chan_Push_mioi_bdwt;
  input r_segment0_ex_ar_chan_Push_mioi_bcwt;
  output r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  input r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_done_sync_vld;
  input r_segment0_ex_ar_chan_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign r_segment0_ex_ar_chan_Push_mioi_bdwt = r_segment0_ex_ar_chan_Push_mioi_oswt
      & master_process_wen;
  assign r_segment0_ex_ar_chan_Push_mioi_biwt = r_segment0_ex_ar_chan_Push_mioi_oswt
      & (~ r_segment0_ex_ar_chan_Push_mioi_bcwt) & r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_done_sync_vld;
  assign r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct
      = master_process_wen & r_segment0_ex_ar_chan_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_dma_cmd_chan_Pop_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_dma_cmd_chan_Pop_mio_wait_dp
    (
  clk, rst_bar, dma_cmd_chan_Pop_mioi_oswt, dma_cmd_chan_Pop_mioi_wen_comp, dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt,
      dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt, dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt,
      dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt, dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt,
      dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt, dma_cmd_chan_Pop_mioi_biwt,
      dma_cmd_chan_Pop_mioi_bdwt, dma_cmd_chan_Pop_mioi_bcwt, dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z,
      dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z, dma_cmd_chan_Pop_mioi_return_total_len_rsc_z,
      dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z, dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z,
      dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z
);
  input clk;
  input rst_bar;
  input dma_cmd_chan_Pop_mioi_oswt;
  output dma_cmd_chan_Pop_mioi_wen_comp;
  output [31:0] dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt;
  output [31:0] dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt;
  output [31:0] dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt;
  output [31:0] dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt;
  output [15:0] dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt;
  output [15:0] dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt;
  input dma_cmd_chan_Pop_mioi_biwt;
  input dma_cmd_chan_Pop_mioi_bdwt;
  output dma_cmd_chan_Pop_mioi_bcwt;
  reg dma_cmd_chan_Pop_mioi_bcwt;
  input [31:0] dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z;
  input [31:0] dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z;
  input [31:0] dma_cmd_chan_Pop_mioi_return_total_len_rsc_z;
  input [31:0] dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z;
  input [15:0] dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z;
  input [15:0] dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z;


  // Interconnect Declarations
  reg [31:0] dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_bfwt;
  reg [31:0] dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_bfwt;
  reg [31:0] dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_bfwt;
  reg [31:0] dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_bfwt;
  reg [15:0] dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_bfwt;
  reg [15:0] dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_cmd_chan_Pop_mioi_wen_comp = (~ dma_cmd_chan_Pop_mioi_oswt) | dma_cmd_chan_Pop_mioi_biwt
      | dma_cmd_chan_Pop_mioi_bcwt;
  assign dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt = MUX_v_32_2_2(dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z,
      dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_bfwt, dma_cmd_chan_Pop_mioi_bcwt);
  assign dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt = MUX_v_32_2_2(dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z,
      dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_bfwt, dma_cmd_chan_Pop_mioi_bcwt);
  assign dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt = MUX_v_32_2_2(dma_cmd_chan_Pop_mioi_return_total_len_rsc_z,
      dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_bfwt, dma_cmd_chan_Pop_mioi_bcwt);
  assign dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt = MUX_v_32_2_2(dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z,
      dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_bfwt, dma_cmd_chan_Pop_mioi_bcwt);
  assign dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt = MUX_v_16_2_2(dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z,
      dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_bfwt, dma_cmd_chan_Pop_mioi_bcwt);
  assign dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt = MUX_v_16_2_2(dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z,
      dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_bfwt, dma_cmd_chan_Pop_mioi_bcwt);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      dma_cmd_chan_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_cmd_chan_Pop_mioi_bcwt <= ~((~(dma_cmd_chan_Pop_mioi_bcwt | dma_cmd_chan_Pop_mioi_biwt))
          | dma_cmd_chan_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_bfwt <= 32'b00000000000000000000000000000000;
      dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_bfwt <= 32'b00000000000000000000000000000000;
      dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_bfwt <= 32'b00000000000000000000000000000000;
      dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_bfwt <= 32'b00000000000000000000000000000000;
      dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_bfwt <= 16'b0000000000000000;
      dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_bfwt <= 16'b0000000000000000;
    end
    else if ( dma_cmd_chan_Pop_mioi_biwt ) begin
      dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_bfwt <= dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z;
      dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_bfwt <= dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z;
      dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_bfwt <= dma_cmd_chan_Pop_mioi_return_total_len_rsc_z;
      dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_bfwt <= dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z;
      dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_bfwt <= dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z;
      dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_bfwt <= dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_dma_cmd_chan_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_dma_cmd_chan_Pop_mio_wait_ctrl
    (
  master_process_wen, dma_cmd_chan_Pop_mioi_oswt, dma_cmd_chan_Pop_mioi_biwt, dma_cmd_chan_Pop_mioi_bdwt,
      dma_cmd_chan_Pop_mioi_bcwt, dma_cmd_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct,
      dma_cmd_chan_Pop_mioi_ccs_ccore_done_sync_vld, dma_cmd_chan_Pop_mioi_oswt_pff
);
  input master_process_wen;
  input dma_cmd_chan_Pop_mioi_oswt;
  output dma_cmd_chan_Pop_mioi_biwt;
  output dma_cmd_chan_Pop_mioi_bdwt;
  input dma_cmd_chan_Pop_mioi_bcwt;
  output dma_cmd_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  input dma_cmd_chan_Pop_mioi_ccs_ccore_done_sync_vld;
  input dma_cmd_chan_Pop_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_cmd_chan_Pop_mioi_bdwt = dma_cmd_chan_Pop_mioi_oswt & master_process_wen;
  assign dma_cmd_chan_Pop_mioi_biwt = dma_cmd_chan_Pop_mioi_oswt & (~ dma_cmd_chan_Pop_mioi_bcwt)
      & dma_cmd_chan_Pop_mioi_ccs_ccore_done_sync_vld;
  assign dma_cmd_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct = master_process_wen
      & dma_cmd_chan_Pop_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_slave_process_fsm
//  FSM Module
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_slave_process_fsm (
  clk, rst_bar, slave_process_wen, fsm_output
);
  input clk;
  input rst_bar;
  input slave_process_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for scatter_gather_dma_slave_process_slave_process_fsm_1
  parameter
    slave_process_rlp_C_0 = 2'd0,
    while_C_0 = 2'd1,
    while_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : scatter_gather_dma_slave_process_slave_process_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = while_C_1;
      end
      while_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = while_C_0;
      end
      // slave_process_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      state_var <= slave_process_rlp_C_0;
    end
    else if ( slave_process_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_staller
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_staller (
  slave_process_wen, w_slave0_aw_Pop_mioi_wen_comp, w_slave0_w_Pop_mioi_wen_comp,
      dma_cmd_chan_Push_mioi_wen_comp, w_slave0_b_Push_mioi_wen_comp
);
  output slave_process_wen;
  input w_slave0_aw_Pop_mioi_wen_comp;
  input w_slave0_w_Pop_mioi_wen_comp;
  input dma_cmd_chan_Push_mioi_wen_comp;
  input w_slave0_b_Push_mioi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign slave_process_wen = w_slave0_aw_Pop_mioi_wen_comp & w_slave0_w_Pop_mioi_wen_comp
      & dma_cmd_chan_Push_mioi_wen_comp & w_slave0_b_Push_mioi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_dp
    (
  clk, rst_bar, w_slave0_b_Push_mioi_oswt, w_slave0_b_Push_mioi_wen_comp, w_slave0_b_Push_mioi_idat_slave_process,
      w_slave0_b_Push_mioi_biwt, w_slave0_b_Push_mioi_bdwt, w_slave0_b_Push_mioi_bcwt,
      w_slave0_b_Push_mioi_idat
);
  input clk;
  input rst_bar;
  input w_slave0_b_Push_mioi_oswt;
  output w_slave0_b_Push_mioi_wen_comp;
  input [1:0] w_slave0_b_Push_mioi_idat_slave_process;
  input w_slave0_b_Push_mioi_biwt;
  input w_slave0_b_Push_mioi_bdwt;
  output w_slave0_b_Push_mioi_bcwt;
  reg w_slave0_b_Push_mioi_bcwt;
  output [1:0] w_slave0_b_Push_mioi_idat;



  // Interconnect Declarations for Component Instantiations 
  assign w_slave0_b_Push_mioi_wen_comp = (~ w_slave0_b_Push_mioi_oswt) | w_slave0_b_Push_mioi_biwt
      | w_slave0_b_Push_mioi_bcwt;
  assign w_slave0_b_Push_mioi_idat = {(w_slave0_b_Push_mioi_idat_slave_process[1])
      , 1'b0};
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_slave0_b_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      w_slave0_b_Push_mioi_bcwt <= ~((~(w_slave0_b_Push_mioi_bcwt | w_slave0_b_Push_mioi_biwt))
          | w_slave0_b_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_ctrl
    (
  slave_process_wen, w_slave0_b_Push_mioi_oswt, w_slave0_b_Push_mioi_biwt, w_slave0_b_Push_mioi_bdwt,
      w_slave0_b_Push_mioi_bcwt, w_slave0_b_Push_mioi_ivld_slave_process_sct, w_slave0_b_Push_mioi_irdy
);
  input slave_process_wen;
  input w_slave0_b_Push_mioi_oswt;
  output w_slave0_b_Push_mioi_biwt;
  output w_slave0_b_Push_mioi_bdwt;
  input w_slave0_b_Push_mioi_bcwt;
  output w_slave0_b_Push_mioi_ivld_slave_process_sct;
  input w_slave0_b_Push_mioi_irdy;


  // Interconnect Declarations
  wire w_slave0_b_Push_mioi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_slave0_b_Push_mioi_bdwt = w_slave0_b_Push_mioi_oswt & slave_process_wen;
  assign w_slave0_b_Push_mioi_biwt = w_slave0_b_Push_mioi_ogwt & w_slave0_b_Push_mioi_irdy;
  assign w_slave0_b_Push_mioi_ogwt = w_slave0_b_Push_mioi_oswt & (~ w_slave0_b_Push_mioi_bcwt);
  assign w_slave0_b_Push_mioi_ivld_slave_process_sct = w_slave0_b_Push_mioi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_dma_cmd_chan_Push_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_dma_cmd_chan_Push_mio_wait_dp
    (
  clk, rst_bar, dma_cmd_chan_Push_mioi_oswt, dma_cmd_chan_Push_mioi_wen_comp, dma_cmd_chan_Push_mioi_biwt,
      dma_cmd_chan_Push_mioi_bdwt, dma_cmd_chan_Push_mioi_bcwt
);
  input clk;
  input rst_bar;
  input dma_cmd_chan_Push_mioi_oswt;
  output dma_cmd_chan_Push_mioi_wen_comp;
  input dma_cmd_chan_Push_mioi_biwt;
  input dma_cmd_chan_Push_mioi_bdwt;
  output dma_cmd_chan_Push_mioi_bcwt;
  reg dma_cmd_chan_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_cmd_chan_Push_mioi_wen_comp = (~ dma_cmd_chan_Push_mioi_oswt) | dma_cmd_chan_Push_mioi_biwt
      | dma_cmd_chan_Push_mioi_bcwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      dma_cmd_chan_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_cmd_chan_Push_mioi_bcwt <= ~((~(dma_cmd_chan_Push_mioi_bcwt | dma_cmd_chan_Push_mioi_biwt))
          | dma_cmd_chan_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_dma_cmd_chan_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_dma_cmd_chan_Push_mio_wait_ctrl
    (
  slave_process_wen, dma_cmd_chan_Push_mioi_oswt, dma_cmd_chan_Push_mioi_biwt, dma_cmd_chan_Push_mioi_bdwt,
      dma_cmd_chan_Push_mioi_bcwt, dma_cmd_chan_Push_mioi_ccs_ccore_start_rsc_dat_slave_process_sct,
      dma_cmd_chan_Push_mioi_ccs_ccore_done_sync_vld, dma_cmd_chan_Push_mioi_oswt_pff
);
  input slave_process_wen;
  input dma_cmd_chan_Push_mioi_oswt;
  output dma_cmd_chan_Push_mioi_biwt;
  output dma_cmd_chan_Push_mioi_bdwt;
  input dma_cmd_chan_Push_mioi_bcwt;
  output dma_cmd_chan_Push_mioi_ccs_ccore_start_rsc_dat_slave_process_sct;
  input dma_cmd_chan_Push_mioi_ccs_ccore_done_sync_vld;
  input dma_cmd_chan_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_cmd_chan_Push_mioi_bdwt = dma_cmd_chan_Push_mioi_oswt & slave_process_wen;
  assign dma_cmd_chan_Push_mioi_biwt = dma_cmd_chan_Push_mioi_oswt & (~ dma_cmd_chan_Push_mioi_bcwt)
      & dma_cmd_chan_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_cmd_chan_Push_mioi_ccs_ccore_start_rsc_dat_slave_process_sct = slave_process_wen
      & dma_cmd_chan_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi_w_slave0_w_Pop_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi_w_slave0_w_Pop_mio_wait_dp
    (
  clk, rst_bar, w_slave0_w_Pop_mioi_oswt, w_slave0_w_Pop_mioi_wen_comp, w_slave0_w_Pop_mioi_idat_mxwt,
      w_slave0_w_Pop_mioi_biwt, w_slave0_w_Pop_mioi_bdwt, w_slave0_w_Pop_mioi_bcwt,
      w_slave0_w_Pop_mioi_idat
);
  input clk;
  input rst_bar;
  input w_slave0_w_Pop_mioi_oswt;
  output w_slave0_w_Pop_mioi_wen_comp;
  output [31:0] w_slave0_w_Pop_mioi_idat_mxwt;
  input w_slave0_w_Pop_mioi_biwt;
  input w_slave0_w_Pop_mioi_bdwt;
  output w_slave0_w_Pop_mioi_bcwt;
  reg w_slave0_w_Pop_mioi_bcwt;
  input [31:0] w_slave0_w_Pop_mioi_idat;


  // Interconnect Declarations
  reg [31:0] w_slave0_w_Pop_mioi_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_slave0_w_Pop_mioi_wen_comp = (~ w_slave0_w_Pop_mioi_oswt) | w_slave0_w_Pop_mioi_biwt
      | w_slave0_w_Pop_mioi_bcwt;
  assign w_slave0_w_Pop_mioi_idat_mxwt = MUX_v_32_2_2(w_slave0_w_Pop_mioi_idat, w_slave0_w_Pop_mioi_idat_bfwt,
      w_slave0_w_Pop_mioi_bcwt);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_slave0_w_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      w_slave0_w_Pop_mioi_bcwt <= ~((~(w_slave0_w_Pop_mioi_bcwt | w_slave0_w_Pop_mioi_biwt))
          | w_slave0_w_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_slave0_w_Pop_mioi_idat_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( w_slave0_w_Pop_mioi_biwt ) begin
      w_slave0_w_Pop_mioi_idat_bfwt <= w_slave0_w_Pop_mioi_idat;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi_w_slave0_w_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi_w_slave0_w_Pop_mio_wait_ctrl
    (
  slave_process_wen, w_slave0_w_Pop_mioi_oswt, w_slave0_w_Pop_mioi_biwt, w_slave0_w_Pop_mioi_bdwt,
      w_slave0_w_Pop_mioi_bcwt, w_slave0_w_Pop_mioi_irdy_slave_process_sct, w_slave0_w_Pop_mioi_ivld
);
  input slave_process_wen;
  input w_slave0_w_Pop_mioi_oswt;
  output w_slave0_w_Pop_mioi_biwt;
  output w_slave0_w_Pop_mioi_bdwt;
  input w_slave0_w_Pop_mioi_bcwt;
  output w_slave0_w_Pop_mioi_irdy_slave_process_sct;
  input w_slave0_w_Pop_mioi_ivld;


  // Interconnect Declarations
  wire w_slave0_w_Pop_mioi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_slave0_w_Pop_mioi_bdwt = w_slave0_w_Pop_mioi_oswt & slave_process_wen;
  assign w_slave0_w_Pop_mioi_biwt = w_slave0_w_Pop_mioi_ogwt & w_slave0_w_Pop_mioi_ivld;
  assign w_slave0_w_Pop_mioi_ogwt = w_slave0_w_Pop_mioi_oswt & (~ w_slave0_w_Pop_mioi_bcwt);
  assign w_slave0_w_Pop_mioi_irdy_slave_process_sct = w_slave0_w_Pop_mioi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi_w_slave0_aw_Pop_mio_wait_dp
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi_w_slave0_aw_Pop_mio_wait_dp
    (
  clk, rst_bar, w_slave0_aw_Pop_mioi_oswt, w_slave0_aw_Pop_mioi_wen_comp, w_slave0_aw_Pop_mioi_idat_mxwt,
      w_slave0_aw_Pop_mioi_biwt, w_slave0_aw_Pop_mioi_bdwt, w_slave0_aw_Pop_mioi_bcwt,
      w_slave0_aw_Pop_mioi_idat
);
  input clk;
  input rst_bar;
  input w_slave0_aw_Pop_mioi_oswt;
  output w_slave0_aw_Pop_mioi_wen_comp;
  output [31:0] w_slave0_aw_Pop_mioi_idat_mxwt;
  input w_slave0_aw_Pop_mioi_biwt;
  input w_slave0_aw_Pop_mioi_bdwt;
  output w_slave0_aw_Pop_mioi_bcwt;
  reg w_slave0_aw_Pop_mioi_bcwt;
  input [31:0] w_slave0_aw_Pop_mioi_idat;


  // Interconnect Declarations
  reg [31:0] w_slave0_aw_Pop_mioi_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_slave0_aw_Pop_mioi_wen_comp = (~ w_slave0_aw_Pop_mioi_oswt) | w_slave0_aw_Pop_mioi_biwt
      | w_slave0_aw_Pop_mioi_bcwt;
  assign w_slave0_aw_Pop_mioi_idat_mxwt = MUX_v_32_2_2(w_slave0_aw_Pop_mioi_idat,
      w_slave0_aw_Pop_mioi_idat_bfwt, w_slave0_aw_Pop_mioi_bcwt);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_slave0_aw_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      w_slave0_aw_Pop_mioi_bcwt <= ~((~(w_slave0_aw_Pop_mioi_bcwt | w_slave0_aw_Pop_mioi_biwt))
          | w_slave0_aw_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_slave0_aw_Pop_mioi_idat_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( w_slave0_aw_Pop_mioi_biwt ) begin
      w_slave0_aw_Pop_mioi_idat_bfwt <= w_slave0_aw_Pop_mioi_idat;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi_w_slave0_aw_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi_w_slave0_aw_Pop_mio_wait_ctrl
    (
  slave_process_wen, w_slave0_aw_Pop_mioi_oswt, w_slave0_aw_Pop_mioi_biwt, w_slave0_aw_Pop_mioi_bdwt,
      w_slave0_aw_Pop_mioi_bcwt, w_slave0_aw_Pop_mioi_irdy_slave_process_sct, w_slave0_aw_Pop_mioi_ivld
);
  input slave_process_wen;
  input w_slave0_aw_Pop_mioi_oswt;
  output w_slave0_aw_Pop_mioi_biwt;
  output w_slave0_aw_Pop_mioi_bdwt;
  input w_slave0_aw_Pop_mioi_bcwt;
  output w_slave0_aw_Pop_mioi_irdy_slave_process_sct;
  input w_slave0_aw_Pop_mioi_ivld;


  // Interconnect Declarations
  wire w_slave0_aw_Pop_mioi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_slave0_aw_Pop_mioi_bdwt = w_slave0_aw_Pop_mioi_oswt & slave_process_wen;
  assign w_slave0_aw_Pop_mioi_biwt = w_slave0_aw_Pop_mioi_ogwt & w_slave0_aw_Pop_mioi_ivld;
  assign w_slave0_aw_Pop_mioi_ogwt = w_slave0_aw_Pop_mioi_oswt & (~ w_slave0_aw_Pop_mioi_bcwt);
  assign w_slave0_aw_Pop_mioi_irdy_slave_process_sct = w_slave0_aw_Pop_mioi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_process_fsm
//  FSM Module
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_process_fsm (
  clk, rst_bar, b_process_wen, fsm_output
);
  input clk;
  input rst_bar;
  input b_process_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_process_fsm_1
  parameter
    b_process_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_process_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // b_process_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      state_var <= b_process_rlp_C_0;
    end
    else if ( b_process_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_staller_2
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_staller_2 (
  clk, rst_bar, b_process_flen_unreg, b_process_wen, b_process_wten, b_in_Pop_mioi_wen_comp,
      last_burst_chan_Pop_mioi_wen_comp, b_chan_Push_mioi_wen_comp
);
  input clk;
  input rst_bar;
  input b_process_flen_unreg;
  output b_process_wen;
  output b_process_wten;
  input b_in_Pop_mioi_wen_comp;
  input last_burst_chan_Pop_mioi_wen_comp;
  input b_chan_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg b_process_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign b_process_wen = b_in_Pop_mioi_wen_comp & last_burst_chan_Pop_mioi_wen_comp
      & b_chan_Push_mioi_wen_comp & (~ b_process_flen_unreg);
  assign b_process_wten = b_process_wten_reg;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      b_process_wten_reg <= 1'b0;
    end
    else begin
      b_process_wten_reg <= ~ b_process_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_b_chan_Push_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_b_chan_Push_mio_wait_dp
    (
  clk, rst_bar, b_chan_Push_mioi_oswt_unreg, b_chan_Push_mioi_bawt, b_chan_Push_mioi_wen_comp,
      b_chan_Push_mioi_biwt, b_chan_Push_mioi_bdwt
);
  input clk;
  input rst_bar;
  input b_chan_Push_mioi_oswt_unreg;
  output b_chan_Push_mioi_bawt;
  output b_chan_Push_mioi_wen_comp;
  input b_chan_Push_mioi_biwt;
  input b_chan_Push_mioi_bdwt;


  // Interconnect Declarations
  reg b_chan_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign b_chan_Push_mioi_bawt = b_chan_Push_mioi_biwt | b_chan_Push_mioi_bcwt;
  assign b_chan_Push_mioi_wen_comp = (~ b_chan_Push_mioi_oswt_unreg) | b_chan_Push_mioi_bawt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      b_chan_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      b_chan_Push_mioi_bcwt <= ~((~(b_chan_Push_mioi_bcwt | b_chan_Push_mioi_biwt))
          | b_chan_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_b_chan_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_b_chan_Push_mio_wait_ctrl
    (
  clk, rst_bar, b_chan_Push_mioi_oswt_unreg, b_process_wen, b_process_wten, b_chan_Push_mioi_iswt0,
      b_chan_Push_mioi_biwt, b_chan_Push_mioi_bdwt, b_chan_Push_mioi_ivld_b_process_sct,
      b_chan_Push_mioi_irdy
);
  input clk;
  input rst_bar;
  input b_chan_Push_mioi_oswt_unreg;
  input b_process_wen;
  input b_process_wten;
  input b_chan_Push_mioi_iswt0;
  output b_chan_Push_mioi_biwt;
  output b_chan_Push_mioi_bdwt;
  output b_chan_Push_mioi_ivld_b_process_sct;
  input b_chan_Push_mioi_irdy;


  // Interconnect Declarations
  wire b_chan_Push_mioi_ogwt;
  reg b_chan_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign b_chan_Push_mioi_bdwt = b_chan_Push_mioi_oswt_unreg & b_process_wen;
  assign b_chan_Push_mioi_biwt = b_chan_Push_mioi_ogwt & b_chan_Push_mioi_irdy;
  assign b_chan_Push_mioi_ogwt = ((~ b_process_wten) & b_chan_Push_mioi_iswt0) |
      b_chan_Push_mioi_icwt;
  assign b_chan_Push_mioi_ivld_b_process_sct = b_chan_Push_mioi_ogwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      b_chan_Push_mioi_icwt <= 1'b0;
    end
    else begin
      b_chan_Push_mioi_icwt <= b_chan_Push_mioi_ogwt & (~ b_chan_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi_last_burst_chan_Pop_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi_last_burst_chan_Pop_mio_wait_dp
    (
  clk, rst_bar, last_burst_chan_Pop_mioi_oswt_unreg, last_burst_chan_Pop_mioi_bawt,
      last_burst_chan_Pop_mioi_wen_comp, last_burst_chan_Pop_mioi_return_rsc_z_mxwt,
      last_burst_chan_Pop_mioi_biwt, last_burst_chan_Pop_mioi_bdwt, last_burst_chan_Pop_mioi_return_rsc_z
);
  input clk;
  input rst_bar;
  input last_burst_chan_Pop_mioi_oswt_unreg;
  output last_burst_chan_Pop_mioi_bawt;
  output last_burst_chan_Pop_mioi_wen_comp;
  output last_burst_chan_Pop_mioi_return_rsc_z_mxwt;
  input last_burst_chan_Pop_mioi_biwt;
  input last_burst_chan_Pop_mioi_bdwt;
  input last_burst_chan_Pop_mioi_return_rsc_z;


  // Interconnect Declarations
  reg last_burst_chan_Pop_mioi_bcwt;
  reg last_burst_chan_Pop_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign last_burst_chan_Pop_mioi_bawt = last_burst_chan_Pop_mioi_biwt | last_burst_chan_Pop_mioi_bcwt;
  assign last_burst_chan_Pop_mioi_wen_comp = (~ last_burst_chan_Pop_mioi_oswt_unreg)
      | last_burst_chan_Pop_mioi_bawt;
  assign last_burst_chan_Pop_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(last_burst_chan_Pop_mioi_return_rsc_z,
      last_burst_chan_Pop_mioi_return_rsc_z_bfwt, last_burst_chan_Pop_mioi_bcwt);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_burst_chan_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      last_burst_chan_Pop_mioi_bcwt <= ~((~(last_burst_chan_Pop_mioi_bcwt | last_burst_chan_Pop_mioi_biwt))
          | last_burst_chan_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_burst_chan_Pop_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( last_burst_chan_Pop_mioi_biwt ) begin
      last_burst_chan_Pop_mioi_return_rsc_z_bfwt <= last_burst_chan_Pop_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi_last_burst_chan_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi_last_burst_chan_Pop_mio_wait_ctrl
    (
  clk, rst_bar, last_burst_chan_Pop_mioi_oswt_unreg, b_process_wen, b_process_wten,
      last_burst_chan_Pop_mioi_iswt0, last_burst_chan_Pop_mioi_biwt, last_burst_chan_Pop_mioi_bdwt,
      last_burst_chan_Pop_mioi_ccs_ccore_start_rsc_dat_b_process_sct, last_burst_chan_Pop_mioi_ccs_ccore_done_sync_vld,
      last_burst_chan_Pop_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  input last_burst_chan_Pop_mioi_oswt_unreg;
  input b_process_wen;
  input b_process_wten;
  input last_burst_chan_Pop_mioi_iswt0;
  output last_burst_chan_Pop_mioi_biwt;
  output last_burst_chan_Pop_mioi_bdwt;
  output last_burst_chan_Pop_mioi_ccs_ccore_start_rsc_dat_b_process_sct;
  input last_burst_chan_Pop_mioi_ccs_ccore_done_sync_vld;
  input last_burst_chan_Pop_mioi_iswt0_pff;


  // Interconnect Declarations
  wire last_burst_chan_Pop_mioi_ogwt;
  reg last_burst_chan_Pop_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign last_burst_chan_Pop_mioi_bdwt = last_burst_chan_Pop_mioi_oswt_unreg & b_process_wen;
  assign last_burst_chan_Pop_mioi_biwt = last_burst_chan_Pop_mioi_ogwt & last_burst_chan_Pop_mioi_ccs_ccore_done_sync_vld;
  assign last_burst_chan_Pop_mioi_ogwt = ((~ b_process_wten) & last_burst_chan_Pop_mioi_iswt0)
      | last_burst_chan_Pop_mioi_icwt;
  assign last_burst_chan_Pop_mioi_ccs_ccore_start_rsc_dat_b_process_sct = b_process_wen
      & last_burst_chan_Pop_mioi_iswt0_pff;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_burst_chan_Pop_mioi_icwt <= 1'b0;
    end
    else begin
      last_burst_chan_Pop_mioi_icwt <= last_burst_chan_Pop_mioi_ogwt & (~ last_burst_chan_Pop_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi_b_in_Pop_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi_b_in_Pop_mio_wait_dp
    (
  clk, rst_bar, b_in_Pop_mioi_oswt_unreg, b_in_Pop_mioi_bawt, b_in_Pop_mioi_wen_comp,
      b_in_Pop_mioi_idat_mxwt, b_in_Pop_mioi_biwt, b_in_Pop_mioi_bdwt, b_in_Pop_mioi_idat
);
  input clk;
  input rst_bar;
  input b_in_Pop_mioi_oswt_unreg;
  output b_in_Pop_mioi_bawt;
  output b_in_Pop_mioi_wen_comp;
  output [5:0] b_in_Pop_mioi_idat_mxwt;
  input b_in_Pop_mioi_biwt;
  input b_in_Pop_mioi_bdwt;
  input [5:0] b_in_Pop_mioi_idat;


  // Interconnect Declarations
  reg b_in_Pop_mioi_bcwt;
  reg [5:0] b_in_Pop_mioi_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign b_in_Pop_mioi_bawt = b_in_Pop_mioi_biwt | b_in_Pop_mioi_bcwt;
  assign b_in_Pop_mioi_wen_comp = (~ b_in_Pop_mioi_oswt_unreg) | b_in_Pop_mioi_bawt;
  assign b_in_Pop_mioi_idat_mxwt = MUX_v_6_2_2(b_in_Pop_mioi_idat, b_in_Pop_mioi_idat_bfwt,
      b_in_Pop_mioi_bcwt);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      b_in_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      b_in_Pop_mioi_bcwt <= ~((~(b_in_Pop_mioi_bcwt | b_in_Pop_mioi_biwt)) | b_in_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      b_in_Pop_mioi_idat_bfwt <= 6'b000000;
    end
    else if ( b_in_Pop_mioi_biwt ) begin
      b_in_Pop_mioi_idat_bfwt <= b_in_Pop_mioi_idat;
    end
  end

  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi_b_in_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi_b_in_Pop_mio_wait_ctrl
    (
  clk, rst_bar, b_in_Pop_mioi_oswt_unreg, b_process_wen, b_process_wten, b_in_Pop_mioi_iswt0,
      b_in_Pop_mioi_biwt, b_in_Pop_mioi_bdwt, b_in_Pop_mioi_irdy_b_process_sct, b_in_Pop_mioi_ivld
);
  input clk;
  input rst_bar;
  input b_in_Pop_mioi_oswt_unreg;
  input b_process_wen;
  input b_process_wten;
  input b_in_Pop_mioi_iswt0;
  output b_in_Pop_mioi_biwt;
  output b_in_Pop_mioi_bdwt;
  output b_in_Pop_mioi_irdy_b_process_sct;
  input b_in_Pop_mioi_ivld;


  // Interconnect Declarations
  wire b_in_Pop_mioi_ogwt;
  reg b_in_Pop_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign b_in_Pop_mioi_bdwt = b_in_Pop_mioi_oswt_unreg & b_process_wen;
  assign b_in_Pop_mioi_biwt = b_in_Pop_mioi_ogwt & b_in_Pop_mioi_ivld;
  assign b_in_Pop_mioi_ogwt = ((~ b_process_wten) & b_in_Pop_mioi_iswt0) | b_in_Pop_mioi_icwt;
  assign b_in_Pop_mioi_irdy_b_process_sct = b_in_Pop_mioi_ogwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      b_in_Pop_mioi_icwt <= 1'b0;
    end
    else begin
      b_in_Pop_mioi_icwt <= b_in_Pop_mioi_ogwt & (~ b_in_Pop_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_process_fsm
//  FSM Module
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_process_fsm (
  clk, rst_bar, w_process_wen, fsm_output
);
  input clk;
  input rst_bar;
  input w_process_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_process_fsm_1
  parameter
    w_process_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_process_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // w_process_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      state_var <= w_process_rlp_C_0;
    end
    else if ( w_process_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_staller_1
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_staller_1 (
  clk, rst_bar, w_process_flen_unreg, w_process_wen, w_process_wten, w_chan_Pop_mioi_wen_comp,
      last_bit_chan_Pop_mioi_wen_comp, w_out_Push_mioi_wen_comp
);
  input clk;
  input rst_bar;
  input w_process_flen_unreg;
  output w_process_wen;
  output w_process_wten;
  input w_chan_Pop_mioi_wen_comp;
  input last_bit_chan_Pop_mioi_wen_comp;
  input w_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg w_process_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign w_process_wen = w_chan_Pop_mioi_wen_comp & last_bit_chan_Pop_mioi_wen_comp
      & w_out_Push_mioi_wen_comp & (~ w_process_flen_unreg);
  assign w_process_wten = w_process_wten_reg;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_process_wten_reg <= 1'b0;
    end
    else begin
      w_process_wten_reg <= ~ w_process_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_w_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_w_out_Push_mio_wait_dp
    (
  clk, rst_bar, w_out_Push_mioi_oswt_unreg, w_out_Push_mioi_bawt, w_out_Push_mioi_wen_comp,
      w_out_Push_mioi_biwt, w_out_Push_mioi_bdwt
);
  input clk;
  input rst_bar;
  input w_out_Push_mioi_oswt_unreg;
  output w_out_Push_mioi_bawt;
  output w_out_Push_mioi_wen_comp;
  input w_out_Push_mioi_biwt;
  input w_out_Push_mioi_bdwt;


  // Interconnect Declarations
  reg w_out_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_out_Push_mioi_bawt = w_out_Push_mioi_biwt | w_out_Push_mioi_bcwt;
  assign w_out_Push_mioi_wen_comp = (~ w_out_Push_mioi_oswt_unreg) | w_out_Push_mioi_bawt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      w_out_Push_mioi_bcwt <= ~((~(w_out_Push_mioi_bcwt | w_out_Push_mioi_biwt))
          | w_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_w_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_w_out_Push_mio_wait_ctrl
    (
  clk, rst_bar, w_out_Push_mioi_oswt_unreg, w_process_wen, w_process_wten, w_out_Push_mioi_iswt0,
      w_out_Push_mioi_biwt, w_out_Push_mioi_bdwt, w_out_Push_mioi_ivld_w_process_sct,
      w_out_Push_mioi_irdy
);
  input clk;
  input rst_bar;
  input w_out_Push_mioi_oswt_unreg;
  input w_process_wen;
  input w_process_wten;
  input w_out_Push_mioi_iswt0;
  output w_out_Push_mioi_biwt;
  output w_out_Push_mioi_bdwt;
  output w_out_Push_mioi_ivld_w_process_sct;
  input w_out_Push_mioi_irdy;


  // Interconnect Declarations
  wire w_out_Push_mioi_ogwt;
  reg w_out_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_out_Push_mioi_bdwt = w_out_Push_mioi_oswt_unreg & w_process_wen;
  assign w_out_Push_mioi_biwt = w_out_Push_mioi_ogwt & w_out_Push_mioi_irdy;
  assign w_out_Push_mioi_ogwt = ((~ w_process_wten) & w_out_Push_mioi_iswt0) | w_out_Push_mioi_icwt;
  assign w_out_Push_mioi_ivld_w_process_sct = w_out_Push_mioi_ogwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_out_Push_mioi_icwt <= 1'b0;
    end
    else begin
      w_out_Push_mioi_icwt <= w_out_Push_mioi_ogwt & (~ w_out_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi_last_bit_chan_Pop_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi_last_bit_chan_Pop_mio_wait_dp
    (
  clk, rst_bar, last_bit_chan_Pop_mioi_oswt_unreg, last_bit_chan_Pop_mioi_bawt, last_bit_chan_Pop_mioi_wen_comp,
      last_bit_chan_Pop_mioi_return_rsc_z_mxwt, last_bit_chan_Pop_mioi_biwt, last_bit_chan_Pop_mioi_bdwt,
      last_bit_chan_Pop_mioi_return_rsc_z
);
  input clk;
  input rst_bar;
  input last_bit_chan_Pop_mioi_oswt_unreg;
  output last_bit_chan_Pop_mioi_bawt;
  output last_bit_chan_Pop_mioi_wen_comp;
  output last_bit_chan_Pop_mioi_return_rsc_z_mxwt;
  input last_bit_chan_Pop_mioi_biwt;
  input last_bit_chan_Pop_mioi_bdwt;
  input last_bit_chan_Pop_mioi_return_rsc_z;


  // Interconnect Declarations
  reg last_bit_chan_Pop_mioi_bcwt;
  reg last_bit_chan_Pop_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign last_bit_chan_Pop_mioi_bawt = last_bit_chan_Pop_mioi_biwt | last_bit_chan_Pop_mioi_bcwt;
  assign last_bit_chan_Pop_mioi_wen_comp = (~ last_bit_chan_Pop_mioi_oswt_unreg)
      | last_bit_chan_Pop_mioi_bawt;
  assign last_bit_chan_Pop_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(last_bit_chan_Pop_mioi_return_rsc_z,
      last_bit_chan_Pop_mioi_return_rsc_z_bfwt, last_bit_chan_Pop_mioi_bcwt);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_bit_chan_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      last_bit_chan_Pop_mioi_bcwt <= ~((~(last_bit_chan_Pop_mioi_bcwt | last_bit_chan_Pop_mioi_biwt))
          | last_bit_chan_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_bit_chan_Pop_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( last_bit_chan_Pop_mioi_biwt ) begin
      last_bit_chan_Pop_mioi_return_rsc_z_bfwt <= last_bit_chan_Pop_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi_last_bit_chan_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi_last_bit_chan_Pop_mio_wait_ctrl
    (
  clk, rst_bar, last_bit_chan_Pop_mioi_oswt_unreg, w_process_wen, w_process_wten,
      last_bit_chan_Pop_mioi_iswt0, last_bit_chan_Pop_mioi_biwt, last_bit_chan_Pop_mioi_bdwt,
      last_bit_chan_Pop_mioi_ccs_ccore_start_rsc_dat_w_process_sct, last_bit_chan_Pop_mioi_ccs_ccore_done_sync_vld,
      last_bit_chan_Pop_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  input last_bit_chan_Pop_mioi_oswt_unreg;
  input w_process_wen;
  input w_process_wten;
  input last_bit_chan_Pop_mioi_iswt0;
  output last_bit_chan_Pop_mioi_biwt;
  output last_bit_chan_Pop_mioi_bdwt;
  output last_bit_chan_Pop_mioi_ccs_ccore_start_rsc_dat_w_process_sct;
  input last_bit_chan_Pop_mioi_ccs_ccore_done_sync_vld;
  input last_bit_chan_Pop_mioi_iswt0_pff;


  // Interconnect Declarations
  wire last_bit_chan_Pop_mioi_ogwt;
  reg last_bit_chan_Pop_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign last_bit_chan_Pop_mioi_bdwt = last_bit_chan_Pop_mioi_oswt_unreg & w_process_wen;
  assign last_bit_chan_Pop_mioi_biwt = last_bit_chan_Pop_mioi_ogwt & last_bit_chan_Pop_mioi_ccs_ccore_done_sync_vld;
  assign last_bit_chan_Pop_mioi_ogwt = ((~ w_process_wten) & last_bit_chan_Pop_mioi_iswt0)
      | last_bit_chan_Pop_mioi_icwt;
  assign last_bit_chan_Pop_mioi_ccs_ccore_start_rsc_dat_w_process_sct = w_process_wen
      & last_bit_chan_Pop_mioi_iswt0_pff;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_bit_chan_Pop_mioi_icwt <= 1'b0;
    end
    else begin
      last_bit_chan_Pop_mioi_icwt <= last_bit_chan_Pop_mioi_ogwt & (~ last_bit_chan_Pop_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi_w_chan_Pop_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi_w_chan_Pop_mio_wait_dp
    (
  clk, rst_bar, w_chan_Pop_mioi_oswt_unreg, w_chan_Pop_mioi_bawt, w_chan_Pop_mioi_wen_comp,
      w_chan_Pop_mioi_idat_mxwt, w_chan_Pop_mioi_biwt, w_chan_Pop_mioi_bdwt, w_chan_Pop_mioi_idat
);
  input clk;
  input rst_bar;
  input w_chan_Pop_mioi_oswt_unreg;
  output w_chan_Pop_mioi_bawt;
  output w_chan_Pop_mioi_wen_comp;
  output [71:0] w_chan_Pop_mioi_idat_mxwt;
  input w_chan_Pop_mioi_biwt;
  input w_chan_Pop_mioi_bdwt;
  input [72:0] w_chan_Pop_mioi_idat;


  // Interconnect Declarations
  reg w_chan_Pop_mioi_bcwt;
  reg [72:0] w_chan_Pop_mioi_idat_bfwt;
  wire [72:0] w_chan_Pop_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  assign w_chan_Pop_mioi_bawt = w_chan_Pop_mioi_biwt | w_chan_Pop_mioi_bcwt;
  assign w_chan_Pop_mioi_wen_comp = (~ w_chan_Pop_mioi_oswt_unreg) | w_chan_Pop_mioi_bawt;
  assign w_chan_Pop_mioi_idat_mxwt_pconst = MUX_v_73_2_2(w_chan_Pop_mioi_idat, w_chan_Pop_mioi_idat_bfwt,
      w_chan_Pop_mioi_bcwt);
  assign w_chan_Pop_mioi_idat_mxwt = {(w_chan_Pop_mioi_idat_mxwt_pconst[72:65]) ,
      (w_chan_Pop_mioi_idat_mxwt_pconst[63:0])};
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_chan_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      w_chan_Pop_mioi_bcwt <= ~((~(w_chan_Pop_mioi_bcwt | w_chan_Pop_mioi_biwt))
          | w_chan_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_chan_Pop_mioi_idat_bfwt <= 73'b0000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( w_chan_Pop_mioi_biwt ) begin
      w_chan_Pop_mioi_idat_bfwt <= w_chan_Pop_mioi_idat;
    end
  end

  function automatic [72:0] MUX_v_73_2_2;
    input [72:0] input_0;
    input [72:0] input_1;
    input  sel;
    reg [72:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_73_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi_w_chan_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi_w_chan_Pop_mio_wait_ctrl
    (
  clk, rst_bar, w_chan_Pop_mioi_oswt_unreg, w_process_wen, w_process_wten, w_chan_Pop_mioi_iswt0,
      w_chan_Pop_mioi_biwt, w_chan_Pop_mioi_bdwt, w_chan_Pop_mioi_irdy_w_process_sct,
      w_chan_Pop_mioi_ivld
);
  input clk;
  input rst_bar;
  input w_chan_Pop_mioi_oswt_unreg;
  input w_process_wen;
  input w_process_wten;
  input w_chan_Pop_mioi_iswt0;
  output w_chan_Pop_mioi_biwt;
  output w_chan_Pop_mioi_bdwt;
  output w_chan_Pop_mioi_irdy_w_process_sct;
  input w_chan_Pop_mioi_ivld;


  // Interconnect Declarations
  wire w_chan_Pop_mioi_ogwt;
  reg w_chan_Pop_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign w_chan_Pop_mioi_bdwt = w_chan_Pop_mioi_oswt_unreg & w_process_wen;
  assign w_chan_Pop_mioi_biwt = w_chan_Pop_mioi_ogwt & w_chan_Pop_mioi_ivld;
  assign w_chan_Pop_mioi_ogwt = ((~ w_process_wten) & w_chan_Pop_mioi_iswt0) | w_chan_Pop_mioi_icwt;
  assign w_chan_Pop_mioi_irdy_w_process_sct = w_chan_Pop_mioi_ogwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_chan_Pop_mioi_icwt <= 1'b0;
    end
    else begin
      w_chan_Pop_mioi_icwt <= w_chan_Pop_mioi_ogwt & (~ w_chan_Pop_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_process_fsm
//  FSM Module
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_process_fsm
    (
  clk, rst_bar, ex_aw_process_wen, fsm_output
);
  input clk;
  input rst_bar;
  input ex_aw_process_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_process_fsm_1
  parameter
    ex_aw_process_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_process_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // ex_aw_process_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      state_var <= ex_aw_process_rlp_C_0;
    end
    else if ( ex_aw_process_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_staller
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_staller (
  clk, rst_bar, ex_aw_process_wen, ex_aw_process_wten, ex_aw_chan_Pop_mioi_wen_comp,
      aw_out_Push_mioi_wen_comp, last_bit_chan_Push_mioi_wen_comp, last_burst_chan_Push_mioi_wen_comp,
      ex_aw_process_flen_unreg
);
  input clk;
  input rst_bar;
  output ex_aw_process_wen;
  output ex_aw_process_wten;
  input ex_aw_chan_Pop_mioi_wen_comp;
  input aw_out_Push_mioi_wen_comp;
  input last_bit_chan_Push_mioi_wen_comp;
  input last_burst_chan_Push_mioi_wen_comp;
  input ex_aw_process_flen_unreg;


  // Interconnect Declarations
  reg ex_aw_process_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign ex_aw_process_wen = ex_aw_chan_Pop_mioi_wen_comp & aw_out_Push_mioi_wen_comp
      & last_bit_chan_Push_mioi_wen_comp & last_burst_chan_Push_mioi_wen_comp & (~
      ex_aw_process_flen_unreg);
  assign ex_aw_process_wten = ex_aw_process_wten_reg;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_aw_process_wten_reg <= 1'b0;
    end
    else begin
      ex_aw_process_wten_reg <= ~ ex_aw_process_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_last_burst_chan_Push_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_last_burst_chan_Push_mio_wait_dp
    (
  clk, rst_bar, last_burst_chan_Push_mioi_oswt_unreg, last_burst_chan_Push_mioi_bawt,
      last_burst_chan_Push_mioi_wen_comp, last_burst_chan_Push_mioi_biwt, last_burst_chan_Push_mioi_bdwt
);
  input clk;
  input rst_bar;
  input last_burst_chan_Push_mioi_oswt_unreg;
  output last_burst_chan_Push_mioi_bawt;
  output last_burst_chan_Push_mioi_wen_comp;
  input last_burst_chan_Push_mioi_biwt;
  input last_burst_chan_Push_mioi_bdwt;


  // Interconnect Declarations
  reg last_burst_chan_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign last_burst_chan_Push_mioi_bawt = last_burst_chan_Push_mioi_biwt | last_burst_chan_Push_mioi_bcwt;
  assign last_burst_chan_Push_mioi_wen_comp = (~ last_burst_chan_Push_mioi_oswt_unreg)
      | last_burst_chan_Push_mioi_bawt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_burst_chan_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      last_burst_chan_Push_mioi_bcwt <= ~((~(last_burst_chan_Push_mioi_bcwt | last_burst_chan_Push_mioi_biwt))
          | last_burst_chan_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_last_burst_chan_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_last_burst_chan_Push_mio_wait_ctrl
    (
  clk, rst_bar, ex_aw_process_wen, ex_aw_process_wten, last_burst_chan_Push_mioi_oswt_unreg,
      last_burst_chan_Push_mioi_iswt0, last_burst_chan_Push_mioi_biwt, last_burst_chan_Push_mioi_bdwt,
      last_burst_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct, last_burst_chan_Push_mioi_ccs_ccore_done_sync_vld,
      last_burst_chan_Push_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  input ex_aw_process_wen;
  input ex_aw_process_wten;
  input last_burst_chan_Push_mioi_oswt_unreg;
  input last_burst_chan_Push_mioi_iswt0;
  output last_burst_chan_Push_mioi_biwt;
  output last_burst_chan_Push_mioi_bdwt;
  output last_burst_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct;
  input last_burst_chan_Push_mioi_ccs_ccore_done_sync_vld;
  input last_burst_chan_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire last_burst_chan_Push_mioi_ogwt;
  reg last_burst_chan_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign last_burst_chan_Push_mioi_bdwt = last_burst_chan_Push_mioi_oswt_unreg &
      ex_aw_process_wen;
  assign last_burst_chan_Push_mioi_biwt = last_burst_chan_Push_mioi_ogwt & last_burst_chan_Push_mioi_ccs_ccore_done_sync_vld;
  assign last_burst_chan_Push_mioi_ogwt = ((~ ex_aw_process_wten) & last_burst_chan_Push_mioi_iswt0)
      | last_burst_chan_Push_mioi_icwt;
  assign last_burst_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct = ex_aw_process_wen
      & last_burst_chan_Push_mioi_iswt0_pff;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_burst_chan_Push_mioi_icwt <= 1'b0;
    end
    else begin
      last_burst_chan_Push_mioi_icwt <= last_burst_chan_Push_mioi_ogwt & (~ last_burst_chan_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_last_bit_chan_Push_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_last_bit_chan_Push_mio_wait_dp
    (
  clk, rst_bar, last_bit_chan_Push_mioi_oswt_unreg, last_bit_chan_Push_mioi_bawt,
      last_bit_chan_Push_mioi_wen_comp, last_bit_chan_Push_mioi_biwt, last_bit_chan_Push_mioi_bdwt
);
  input clk;
  input rst_bar;
  input last_bit_chan_Push_mioi_oswt_unreg;
  output last_bit_chan_Push_mioi_bawt;
  output last_bit_chan_Push_mioi_wen_comp;
  input last_bit_chan_Push_mioi_biwt;
  input last_bit_chan_Push_mioi_bdwt;


  // Interconnect Declarations
  reg last_bit_chan_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign last_bit_chan_Push_mioi_bawt = last_bit_chan_Push_mioi_biwt | last_bit_chan_Push_mioi_bcwt;
  assign last_bit_chan_Push_mioi_wen_comp = (~ last_bit_chan_Push_mioi_oswt_unreg)
      | last_bit_chan_Push_mioi_bawt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_bit_chan_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      last_bit_chan_Push_mioi_bcwt <= ~((~(last_bit_chan_Push_mioi_bcwt | last_bit_chan_Push_mioi_biwt))
          | last_bit_chan_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_last_bit_chan_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_last_bit_chan_Push_mio_wait_ctrl
    (
  clk, rst_bar, ex_aw_process_wen, ex_aw_process_wten, last_bit_chan_Push_mioi_oswt_unreg,
      last_bit_chan_Push_mioi_iswt0, last_bit_chan_Push_mioi_biwt, last_bit_chan_Push_mioi_bdwt,
      last_bit_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct, last_bit_chan_Push_mioi_ccs_ccore_done_sync_vld,
      last_bit_chan_Push_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  input ex_aw_process_wen;
  input ex_aw_process_wten;
  input last_bit_chan_Push_mioi_oswt_unreg;
  input last_bit_chan_Push_mioi_iswt0;
  output last_bit_chan_Push_mioi_biwt;
  output last_bit_chan_Push_mioi_bdwt;
  output last_bit_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct;
  input last_bit_chan_Push_mioi_ccs_ccore_done_sync_vld;
  input last_bit_chan_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire last_bit_chan_Push_mioi_ogwt;
  reg last_bit_chan_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign last_bit_chan_Push_mioi_bdwt = last_bit_chan_Push_mioi_oswt_unreg & ex_aw_process_wen;
  assign last_bit_chan_Push_mioi_biwt = last_bit_chan_Push_mioi_ogwt & last_bit_chan_Push_mioi_ccs_ccore_done_sync_vld;
  assign last_bit_chan_Push_mioi_ogwt = ((~ ex_aw_process_wten) & last_bit_chan_Push_mioi_iswt0)
      | last_bit_chan_Push_mioi_icwt;
  assign last_bit_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct = ex_aw_process_wen
      & last_bit_chan_Push_mioi_iswt0_pff;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      last_bit_chan_Push_mioi_icwt <= 1'b0;
    end
    else begin
      last_bit_chan_Push_mioi_icwt <= last_bit_chan_Push_mioi_ogwt & (~ last_bit_chan_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_aw_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_aw_out_Push_mio_wait_dp
    (
  clk, rst_bar, aw_out_Push_mioi_oswt_unreg, aw_out_Push_mioi_bawt, aw_out_Push_mioi_wen_comp,
      aw_out_Push_mioi_biwt, aw_out_Push_mioi_bdwt
);
  input clk;
  input rst_bar;
  input aw_out_Push_mioi_oswt_unreg;
  output aw_out_Push_mioi_bawt;
  output aw_out_Push_mioi_wen_comp;
  input aw_out_Push_mioi_biwt;
  input aw_out_Push_mioi_bdwt;


  // Interconnect Declarations
  reg aw_out_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign aw_out_Push_mioi_bawt = aw_out_Push_mioi_biwt | aw_out_Push_mioi_bcwt;
  assign aw_out_Push_mioi_wen_comp = (~ aw_out_Push_mioi_oswt_unreg) | aw_out_Push_mioi_bawt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      aw_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      aw_out_Push_mioi_bcwt <= ~((~(aw_out_Push_mioi_bcwt | aw_out_Push_mioi_biwt))
          | aw_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_aw_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_aw_out_Push_mio_wait_ctrl
    (
  clk, rst_bar, ex_aw_process_wen, ex_aw_process_wten, aw_out_Push_mioi_oswt_unreg,
      aw_out_Push_mioi_iswt0, aw_out_Push_mioi_biwt, aw_out_Push_mioi_bdwt, aw_out_Push_mioi_ivld_ex_aw_process_sct,
      aw_out_Push_mioi_irdy
);
  input clk;
  input rst_bar;
  input ex_aw_process_wen;
  input ex_aw_process_wten;
  input aw_out_Push_mioi_oswt_unreg;
  input aw_out_Push_mioi_iswt0;
  output aw_out_Push_mioi_biwt;
  output aw_out_Push_mioi_bdwt;
  output aw_out_Push_mioi_ivld_ex_aw_process_sct;
  input aw_out_Push_mioi_irdy;


  // Interconnect Declarations
  wire aw_out_Push_mioi_ogwt;
  reg aw_out_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign aw_out_Push_mioi_bdwt = aw_out_Push_mioi_oswt_unreg & ex_aw_process_wen;
  assign aw_out_Push_mioi_biwt = aw_out_Push_mioi_ogwt & aw_out_Push_mioi_irdy;
  assign aw_out_Push_mioi_ogwt = ((~ ex_aw_process_wten) & aw_out_Push_mioi_iswt0)
      | aw_out_Push_mioi_icwt;
  assign aw_out_Push_mioi_ivld_ex_aw_process_sct = aw_out_Push_mioi_ogwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      aw_out_Push_mioi_icwt <= 1'b0;
    end
    else begin
      aw_out_Push_mioi_icwt <= aw_out_Push_mioi_ogwt & (~ aw_out_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_ex_aw_chan_Pop_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_ex_aw_chan_Pop_mio_wait_dp
    (
  clk, rst_bar, ex_aw_chan_Pop_mioi_oswt_unreg, ex_aw_chan_Pop_mioi_bawt, ex_aw_chan_Pop_mioi_wen_comp,
      ex_aw_chan_Pop_mioi_idat_mxwt, ex_aw_chan_Pop_mioi_biwt, ex_aw_chan_Pop_mioi_bdwt,
      ex_aw_chan_Pop_mioi_idat
);
  input clk;
  input rst_bar;
  input ex_aw_chan_Pop_mioi_oswt_unreg;
  output ex_aw_chan_Pop_mioi_bawt;
  output ex_aw_chan_Pop_mioi_wen_comp;
  output [67:0] ex_aw_chan_Pop_mioi_idat_mxwt;
  input ex_aw_chan_Pop_mioi_biwt;
  input ex_aw_chan_Pop_mioi_bdwt;
  input [75:0] ex_aw_chan_Pop_mioi_idat;


  // Interconnect Declarations
  reg ex_aw_chan_Pop_mioi_bcwt;
  reg [75:0] ex_aw_chan_Pop_mioi_idat_bfwt;
  wire [75:0] ex_aw_chan_Pop_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  assign ex_aw_chan_Pop_mioi_bawt = ex_aw_chan_Pop_mioi_biwt | ex_aw_chan_Pop_mioi_bcwt;
  assign ex_aw_chan_Pop_mioi_wen_comp = (~ ex_aw_chan_Pop_mioi_oswt_unreg) | ex_aw_chan_Pop_mioi_bawt;
  assign ex_aw_chan_Pop_mioi_idat_mxwt_pconst = MUX_v_76_2_2(ex_aw_chan_Pop_mioi_idat,
      ex_aw_chan_Pop_mioi_idat_bfwt, ex_aw_chan_Pop_mioi_bcwt);
  assign ex_aw_chan_Pop_mioi_idat_mxwt = {(ex_aw_chan_Pop_mioi_idat_mxwt_pconst[75:44])
      , (ex_aw_chan_Pop_mioi_idat_mxwt_pconst[35:0])};
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_aw_chan_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      ex_aw_chan_Pop_mioi_bcwt <= ~((~(ex_aw_chan_Pop_mioi_bcwt | ex_aw_chan_Pop_mioi_biwt))
          | ex_aw_chan_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_aw_chan_Pop_mioi_idat_bfwt <= 76'b0000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ex_aw_chan_Pop_mioi_biwt ) begin
      ex_aw_chan_Pop_mioi_idat_bfwt <= ex_aw_chan_Pop_mioi_idat;
    end
  end

  function automatic [75:0] MUX_v_76_2_2;
    input [75:0] input_0;
    input [75:0] input_1;
    input  sel;
    reg [75:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_76_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_ex_aw_chan_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_ex_aw_chan_Pop_mio_wait_ctrl
    (
  clk, rst_bar, ex_aw_process_wen, ex_aw_process_wten, ex_aw_chan_Pop_mioi_oswt_unreg,
      ex_aw_chan_Pop_mioi_iswt0, ex_aw_chan_Pop_mioi_biwt, ex_aw_chan_Pop_mioi_bdwt,
      ex_aw_chan_Pop_mioi_irdy_ex_aw_process_sct, ex_aw_chan_Pop_mioi_ivld
);
  input clk;
  input rst_bar;
  input ex_aw_process_wen;
  input ex_aw_process_wten;
  input ex_aw_chan_Pop_mioi_oswt_unreg;
  input ex_aw_chan_Pop_mioi_iswt0;
  output ex_aw_chan_Pop_mioi_biwt;
  output ex_aw_chan_Pop_mioi_bdwt;
  output ex_aw_chan_Pop_mioi_irdy_ex_aw_process_sct;
  input ex_aw_chan_Pop_mioi_ivld;


  // Interconnect Declarations
  wire ex_aw_chan_Pop_mioi_ogwt;
  reg ex_aw_chan_Pop_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign ex_aw_chan_Pop_mioi_bdwt = ex_aw_chan_Pop_mioi_oswt_unreg & ex_aw_process_wen;
  assign ex_aw_chan_Pop_mioi_biwt = ex_aw_chan_Pop_mioi_ogwt & ex_aw_chan_Pop_mioi_ivld;
  assign ex_aw_chan_Pop_mioi_ogwt = ((~ ex_aw_process_wten) & ex_aw_chan_Pop_mioi_iswt0)
      | ex_aw_chan_Pop_mioi_icwt;
  assign ex_aw_chan_Pop_mioi_irdy_ex_aw_process_sct = ex_aw_chan_Pop_mioi_ogwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_aw_chan_Pop_mioi_icwt <= 1'b0;
    end
    else begin
      ex_aw_chan_Pop_mioi_icwt <= ex_aw_chan_Pop_mioi_ogwt & (~ ex_aw_chan_Pop_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_process_fsm
//  FSM Module
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_process_fsm
    (
  clk, rst_bar, ex_ar_process_wen, fsm_output
);
  input clk;
  input rst_bar;
  input ex_ar_process_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_process_fsm_1
  parameter
    ex_ar_process_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_process_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // ex_ar_process_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      state_var <= ex_ar_process_rlp_C_0;
    end
    else if ( ex_ar_process_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_staller
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_staller (
  clk, rst_bar, ex_ar_process_wen, ex_ar_process_wten, ex_ar_chan_Pop_mioi_wen_comp,
      ar_out_Push_mioi_wen_comp, ex_ar_process_flen_unreg
);
  input clk;
  input rst_bar;
  output ex_ar_process_wen;
  output ex_ar_process_wten;
  reg ex_ar_process_wten;
  input ex_ar_chan_Pop_mioi_wen_comp;
  input ar_out_Push_mioi_wen_comp;
  input ex_ar_process_flen_unreg;



  // Interconnect Declarations for Component Instantiations 
  assign ex_ar_process_wen = ex_ar_chan_Pop_mioi_wen_comp & ar_out_Push_mioi_wen_comp
      & (~ ex_ar_process_flen_unreg);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_ar_process_wten <= 1'b0;
    end
    else begin
      ex_ar_process_wten <= ~ ex_ar_process_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_ar_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_ar_out_Push_mio_wait_dp
    (
  clk, rst_bar, ar_out_Push_mioi_oswt_unreg, ar_out_Push_mioi_bawt, ar_out_Push_mioi_wen_comp,
      ar_out_Push_mioi_biwt, ar_out_Push_mioi_bdwt
);
  input clk;
  input rst_bar;
  input ar_out_Push_mioi_oswt_unreg;
  output ar_out_Push_mioi_bawt;
  output ar_out_Push_mioi_wen_comp;
  input ar_out_Push_mioi_biwt;
  input ar_out_Push_mioi_bdwt;


  // Interconnect Declarations
  reg ar_out_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign ar_out_Push_mioi_bawt = ar_out_Push_mioi_biwt | ar_out_Push_mioi_bcwt;
  assign ar_out_Push_mioi_wen_comp = (~ ar_out_Push_mioi_oswt_unreg) | ar_out_Push_mioi_bawt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ar_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      ar_out_Push_mioi_bcwt <= ~((~(ar_out_Push_mioi_bcwt | ar_out_Push_mioi_biwt))
          | ar_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_ar_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_ar_out_Push_mio_wait_ctrl
    (
  clk, rst_bar, ex_ar_process_wen, ex_ar_process_wten, ar_out_Push_mioi_oswt_unreg,
      ar_out_Push_mioi_iswt0, ar_out_Push_mioi_biwt, ar_out_Push_mioi_bdwt, ar_out_Push_mioi_ivld_ex_ar_process_sct,
      ar_out_Push_mioi_irdy
);
  input clk;
  input rst_bar;
  input ex_ar_process_wen;
  input ex_ar_process_wten;
  input ar_out_Push_mioi_oswt_unreg;
  input ar_out_Push_mioi_iswt0;
  output ar_out_Push_mioi_biwt;
  output ar_out_Push_mioi_bdwt;
  output ar_out_Push_mioi_ivld_ex_ar_process_sct;
  input ar_out_Push_mioi_irdy;


  // Interconnect Declarations
  wire ar_out_Push_mioi_ogwt;
  reg ar_out_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign ar_out_Push_mioi_bdwt = ar_out_Push_mioi_oswt_unreg & ex_ar_process_wen;
  assign ar_out_Push_mioi_biwt = ar_out_Push_mioi_ogwt & ar_out_Push_mioi_irdy;
  assign ar_out_Push_mioi_ogwt = ((~ ex_ar_process_wten) & ar_out_Push_mioi_iswt0)
      | ar_out_Push_mioi_icwt;
  assign ar_out_Push_mioi_ivld_ex_ar_process_sct = ar_out_Push_mioi_ogwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ar_out_Push_mioi_icwt <= 1'b0;
    end
    else begin
      ar_out_Push_mioi_icwt <= ar_out_Push_mioi_ogwt & (~ ar_out_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_ex_ar_chan_Pop_mio_wait_dp
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_ex_ar_chan_Pop_mio_wait_dp
    (
  clk, rst_bar, ex_ar_chan_Pop_mioi_oswt_unreg, ex_ar_chan_Pop_mioi_bawt, ex_ar_chan_Pop_mioi_wen_comp,
      ex_ar_chan_Pop_mioi_idat_mxwt, ex_ar_chan_Pop_mioi_biwt, ex_ar_chan_Pop_mioi_bdwt,
      ex_ar_chan_Pop_mioi_idat
);
  input clk;
  input rst_bar;
  input ex_ar_chan_Pop_mioi_oswt_unreg;
  output ex_ar_chan_Pop_mioi_bawt;
  output ex_ar_chan_Pop_mioi_wen_comp;
  output [67:0] ex_ar_chan_Pop_mioi_idat_mxwt;
  input ex_ar_chan_Pop_mioi_biwt;
  input ex_ar_chan_Pop_mioi_bdwt;
  input [75:0] ex_ar_chan_Pop_mioi_idat;


  // Interconnect Declarations
  reg ex_ar_chan_Pop_mioi_bcwt;
  reg [75:0] ex_ar_chan_Pop_mioi_idat_bfwt;
  wire [75:0] ex_ar_chan_Pop_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  assign ex_ar_chan_Pop_mioi_bawt = ex_ar_chan_Pop_mioi_biwt | ex_ar_chan_Pop_mioi_bcwt;
  assign ex_ar_chan_Pop_mioi_wen_comp = (~ ex_ar_chan_Pop_mioi_oswt_unreg) | ex_ar_chan_Pop_mioi_bawt;
  assign ex_ar_chan_Pop_mioi_idat_mxwt_pconst = MUX_v_76_2_2(ex_ar_chan_Pop_mioi_idat,
      ex_ar_chan_Pop_mioi_idat_bfwt, ex_ar_chan_Pop_mioi_bcwt);
  assign ex_ar_chan_Pop_mioi_idat_mxwt = {(ex_ar_chan_Pop_mioi_idat_mxwt_pconst[75:44])
      , (ex_ar_chan_Pop_mioi_idat_mxwt_pconst[35:0])};
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_ar_chan_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      ex_ar_chan_Pop_mioi_bcwt <= ~((~(ex_ar_chan_Pop_mioi_bcwt | ex_ar_chan_Pop_mioi_biwt))
          | ex_ar_chan_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_ar_chan_Pop_mioi_idat_bfwt <= 76'b0000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ex_ar_chan_Pop_mioi_biwt ) begin
      ex_ar_chan_Pop_mioi_idat_bfwt <= ex_ar_chan_Pop_mioi_idat;
    end
  end

  function automatic [75:0] MUX_v_76_2_2;
    input [75:0] input_0;
    input [75:0] input_1;
    input  sel;
    reg [75:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_76_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_ex_ar_chan_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_ex_ar_chan_Pop_mio_wait_ctrl
    (
  clk, rst_bar, ex_ar_process_wen, ex_ar_process_wten, ex_ar_chan_Pop_mioi_oswt_unreg,
      ex_ar_chan_Pop_mioi_iswt0, ex_ar_chan_Pop_mioi_biwt, ex_ar_chan_Pop_mioi_bdwt,
      ex_ar_chan_Pop_mioi_irdy_ex_ar_process_sct, ex_ar_chan_Pop_mioi_ivld
);
  input clk;
  input rst_bar;
  input ex_ar_process_wen;
  input ex_ar_process_wten;
  input ex_ar_chan_Pop_mioi_oswt_unreg;
  input ex_ar_chan_Pop_mioi_iswt0;
  output ex_ar_chan_Pop_mioi_biwt;
  output ex_ar_chan_Pop_mioi_bdwt;
  output ex_ar_chan_Pop_mioi_irdy_ex_ar_process_sct;
  input ex_ar_chan_Pop_mioi_ivld;


  // Interconnect Declarations
  wire ex_ar_chan_Pop_mioi_ogwt;
  reg ex_ar_chan_Pop_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign ex_ar_chan_Pop_mioi_bdwt = ex_ar_chan_Pop_mioi_oswt_unreg & ex_ar_process_wen;
  assign ex_ar_chan_Pop_mioi_biwt = ex_ar_chan_Pop_mioi_ogwt & ex_ar_chan_Pop_mioi_ivld;
  assign ex_ar_chan_Pop_mioi_ogwt = ((~ ex_ar_process_wten) & ex_ar_chan_Pop_mioi_iswt0)
      | ex_ar_chan_Pop_mioi_icwt;
  assign ex_ar_chan_Pop_mioi_irdy_ex_ar_process_sct = ex_ar_chan_Pop_mioi_ogwt;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_ar_chan_Pop_mioi_icwt <= 1'b0;
    end
    else begin
      ex_ar_chan_Pop_mioi_icwt <= ex_ar_chan_Pop_mioi_ogwt & (~ ex_ar_chan_Pop_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_dma_done_Push_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_dma_done_Push_mioi (
  clk, rst_bar, dma_done_vld, dma_done_rdy, dma_done_dat, master_process_wen, dma_done_Push_mioi_oswt,
      dma_done_Push_mioi_wen_comp, dma_done_Push_mioi_idat_master_process
);
  input clk;
  input rst_bar;
  output dma_done_vld;
  input dma_done_rdy;
  output dma_done_dat;
  input master_process_wen;
  input dma_done_Push_mioi_oswt;
  output dma_done_Push_mioi_wen_comp;
  input dma_done_Push_mioi_idat_master_process;


  // Interconnect Declarations
  wire dma_done_Push_mioi_biwt;
  wire dma_done_Push_mioi_bdwt;
  wire dma_done_Push_mioi_bcwt;
  wire dma_done_Push_mioi_idat_master_process_sct;
  wire dma_done_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_out_wait_v1 #(.width(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) dma_done_Push_mioi (
      .vld(dma_done_vld),
      .rdy(dma_done_rdy),
      .dat(dma_done_dat),
      .idat(dma_done_Push_mioi_idat_master_process),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1),
      .ivld(dma_done_Push_mioi_idat_master_process_sct),
      .irdy(dma_done_Push_mioi_irdy)
    );
  scatter_gather_dma_master_process_dma_done_Push_mioi_dma_done_Push_mio_wait_ctrl
      scatter_gather_dma_master_process_dma_done_Push_mioi_dma_done_Push_mio_wait_ctrl_inst
      (
      .master_process_wen(master_process_wen),
      .dma_done_Push_mioi_oswt(dma_done_Push_mioi_oswt),
      .dma_done_Push_mioi_biwt(dma_done_Push_mioi_biwt),
      .dma_done_Push_mioi_bdwt(dma_done_Push_mioi_bdwt),
      .dma_done_Push_mioi_bcwt(dma_done_Push_mioi_bcwt),
      .dma_done_Push_mioi_idat_master_process_sct(dma_done_Push_mioi_idat_master_process_sct),
      .dma_done_Push_mioi_irdy(dma_done_Push_mioi_irdy)
    );
  scatter_gather_dma_master_process_dma_done_Push_mioi_dma_done_Push_mio_wait_dp
      scatter_gather_dma_master_process_dma_done_Push_mioi_dma_done_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .dma_done_Push_mioi_oswt(dma_done_Push_mioi_oswt),
      .dma_done_Push_mioi_wen_comp(dma_done_Push_mioi_wen_comp),
      .dma_done_Push_mioi_biwt(dma_done_Push_mioi_biwt),
      .dma_done_Push_mioi_bdwt(dma_done_Push_mioi_bdwt),
      .dma_done_Push_mioi_bcwt(dma_done_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi (
  clk, rst_bar, w_segment0_b_chan_vld, w_segment0_b_chan_rdy, w_segment0_b_chan_dat,
      master_process_wen, w_segment0_b_chan_Pop_mioi_oswt, w_segment0_b_chan_Pop_mioi_wen_comp,
      w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt, w_segment0_b_chan_Pop_mioi_oswt_pff
);
  input clk;
  input rst_bar;
  input w_segment0_b_chan_vld;
  output w_segment0_b_chan_rdy;
  input [5:0] w_segment0_b_chan_dat;
  input master_process_wen;
  input w_segment0_b_chan_Pop_mioi_oswt;
  output w_segment0_b_chan_Pop_mioi_wen_comp;
  output [1:0] w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt;
  input w_segment0_b_chan_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire w_segment0_b_chan_Pop_mioi_biwt;
  wire w_segment0_b_chan_Pop_mioi_bdwt;
  wire w_segment0_b_chan_Pop_mioi_bcwt;
  wire [3:0] w_segment0_b_chan_Pop_mioi_return_id_rsc_z;
  wire [1:0] w_segment0_b_chan_Pop_mioi_return_resp_rsc_z;
  wire w_segment0_b_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  wire w_segment0_b_chan_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_axi_axi4_axi_cfg_standard_WRespPayload_Connections_SYN_PORT_Pop
      w_segment0_b_chan_Pop_mioi (
      .this_vld(w_segment0_b_chan_vld),
      .this_rdy(w_segment0_b_chan_rdy),
      .this_dat(w_segment0_b_chan_dat),
      .return_id_rsc_z(w_segment0_b_chan_Pop_mioi_return_id_rsc_z),
      .return_resp_rsc_z(w_segment0_b_chan_Pop_mioi_return_resp_rsc_z),
      .ccs_ccore_start_rsc_dat(w_segment0_b_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .ccs_ccore_done_sync_vld(w_segment0_b_chan_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi_w_segment0_b_chan_Pop_mio_wait_ctrl
      scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi_w_segment0_b_chan_Pop_mio_wait_ctrl_inst
      (
      .master_process_wen(master_process_wen),
      .w_segment0_b_chan_Pop_mioi_oswt(w_segment0_b_chan_Pop_mioi_oswt),
      .w_segment0_b_chan_Pop_mioi_biwt(w_segment0_b_chan_Pop_mioi_biwt),
      .w_segment0_b_chan_Pop_mioi_bdwt(w_segment0_b_chan_Pop_mioi_bdwt),
      .w_segment0_b_chan_Pop_mioi_bcwt(w_segment0_b_chan_Pop_mioi_bcwt),
      .w_segment0_b_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct(w_segment0_b_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .w_segment0_b_chan_Pop_mioi_ccs_ccore_done_sync_vld(w_segment0_b_chan_Pop_mioi_ccs_ccore_done_sync_vld),
      .w_segment0_b_chan_Pop_mioi_oswt_pff(w_segment0_b_chan_Pop_mioi_oswt_pff)
    );
  scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi_w_segment0_b_chan_Pop_mio_wait_dp
      scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi_w_segment0_b_chan_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_segment0_b_chan_Pop_mioi_oswt(w_segment0_b_chan_Pop_mioi_oswt),
      .w_segment0_b_chan_Pop_mioi_wen_comp(w_segment0_b_chan_Pop_mioi_wen_comp),
      .w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt(w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt),
      .w_segment0_b_chan_Pop_mioi_biwt(w_segment0_b_chan_Pop_mioi_biwt),
      .w_segment0_b_chan_Pop_mioi_bdwt(w_segment0_b_chan_Pop_mioi_bdwt),
      .w_segment0_b_chan_Pop_mioi_bcwt(w_segment0_b_chan_Pop_mioi_bcwt),
      .w_segment0_b_chan_Pop_mioi_return_resp_rsc_z(w_segment0_b_chan_Pop_mioi_return_resp_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi (
  clk, rst_bar, w_segment0_w_chan_vld, w_segment0_w_chan_rdy, w_segment0_w_chan_dat,
      w_segment0_w_chan_Push_mioi_oswt_unreg, master_process_wen, master_process_wten,
      w_segment0_w_chan_Push_mioi_bawt, w_segment0_w_chan_Push_mioi_iswt0, w_segment0_w_chan_Push_mioi_wen_comp,
      w_segment0_w_chan_Push_mioi_m_data_rsc_dat, w_segment0_w_chan_Push_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  output w_segment0_w_chan_vld;
  input w_segment0_w_chan_rdy;
  output [72:0] w_segment0_w_chan_dat;
  input w_segment0_w_chan_Push_mioi_oswt_unreg;
  input master_process_wen;
  input master_process_wten;
  output w_segment0_w_chan_Push_mioi_bawt;
  input w_segment0_w_chan_Push_mioi_iswt0;
  output w_segment0_w_chan_Push_mioi_wen_comp;
  input [63:0] w_segment0_w_chan_Push_mioi_m_data_rsc_dat;
  input w_segment0_w_chan_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire w_segment0_w_chan_Push_mioi_biwt;
  wire w_segment0_w_chan_Push_mioi_bdwt;
  wire w_segment0_w_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  wire w_segment0_w_chan_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_Push
      w_segment0_w_chan_Push_mioi (
      .this_vld(w_segment0_w_chan_vld),
      .this_rdy(w_segment0_w_chan_rdy),
      .this_dat(w_segment0_w_chan_dat),
      .m_data_rsc_dat(w_segment0_w_chan_Push_mioi_m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(w_segment0_w_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .ccs_ccore_done_sync_vld(w_segment0_w_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_w_segment0_w_chan_Push_mio_wait_ctrl
      scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_w_segment0_w_chan_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_segment0_w_chan_Push_mioi_oswt_unreg(w_segment0_w_chan_Push_mioi_oswt_unreg),
      .master_process_wen(master_process_wen),
      .master_process_wten(master_process_wten),
      .w_segment0_w_chan_Push_mioi_iswt0(w_segment0_w_chan_Push_mioi_iswt0),
      .w_segment0_w_chan_Push_mioi_biwt(w_segment0_w_chan_Push_mioi_biwt),
      .w_segment0_w_chan_Push_mioi_bdwt(w_segment0_w_chan_Push_mioi_bdwt),
      .w_segment0_w_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct(w_segment0_w_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .w_segment0_w_chan_Push_mioi_ccs_ccore_done_sync_vld(w_segment0_w_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .w_segment0_w_chan_Push_mioi_iswt0_pff(w_segment0_w_chan_Push_mioi_iswt0_pff)
    );
  scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_w_segment0_w_chan_Push_mio_wait_dp
      scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_w_segment0_w_chan_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_segment0_w_chan_Push_mioi_oswt_unreg(w_segment0_w_chan_Push_mioi_oswt_unreg),
      .w_segment0_w_chan_Push_mioi_bawt(w_segment0_w_chan_Push_mioi_bawt),
      .w_segment0_w_chan_Push_mioi_wen_comp(w_segment0_w_chan_Push_mioi_wen_comp),
      .w_segment0_w_chan_Push_mioi_biwt(w_segment0_w_chan_Push_mioi_biwt),
      .w_segment0_w_chan_Push_mioi_bdwt(w_segment0_w_chan_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_r_master0_r_Pop_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_r_master0_r_Pop_mioi (
  clk, rst_bar, r_master0_r_vld, r_master0_r_rdy, r_master0_r_dat, r_master0_r_Pop_mioi_oswt_unreg,
      master_process_wen, master_process_wten, r_master0_r_Pop_mioi_bawt, r_master0_r_Pop_mioi_iswt0,
      r_master0_r_Pop_mioi_wen_comp, r_master0_r_Pop_mioi_idat_mxwt
);
  input clk;
  input rst_bar;
  input r_master0_r_vld;
  output r_master0_r_rdy;
  input [70:0] r_master0_r_dat;
  input r_master0_r_Pop_mioi_oswt_unreg;
  input master_process_wen;
  input master_process_wten;
  output r_master0_r_Pop_mioi_bawt;
  input r_master0_r_Pop_mioi_iswt0;
  output r_master0_r_Pop_mioi_wen_comp;
  output [63:0] r_master0_r_Pop_mioi_idat_mxwt;


  // Interconnect Declarations
  wire r_master0_r_Pop_mioi_biwt;
  wire r_master0_r_Pop_mioi_bdwt;
  wire [70:0] r_master0_r_Pop_mioi_idat;
  wire r_master0_r_Pop_mioi_irdy_master_process_sct;
  wire r_master0_r_Pop_mioi_ivld;
  wire [63:0] r_master0_r_Pop_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_in_wait_v1 #(.width(32'sd71),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) r_master0_r_Pop_mioi (
      .vld(r_master0_r_vld),
      .rdy(r_master0_r_rdy),
      .dat(r_master0_r_dat),
      .idat(r_master0_r_Pop_mioi_idat),
      .irdy(r_master0_r_Pop_mioi_irdy_master_process_sct),
      .ivld(r_master0_r_Pop_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1)
    );
  scatter_gather_dma_master_process_r_master0_r_Pop_mioi_r_master0_r_Pop_mio_wait_ctrl
      scatter_gather_dma_master_process_r_master0_r_Pop_mioi_r_master0_r_Pop_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .r_master0_r_Pop_mioi_oswt_unreg(r_master0_r_Pop_mioi_oswt_unreg),
      .master_process_wen(master_process_wen),
      .master_process_wten(master_process_wten),
      .r_master0_r_Pop_mioi_iswt0(r_master0_r_Pop_mioi_iswt0),
      .r_master0_r_Pop_mioi_biwt(r_master0_r_Pop_mioi_biwt),
      .r_master0_r_Pop_mioi_bdwt(r_master0_r_Pop_mioi_bdwt),
      .r_master0_r_Pop_mioi_irdy_master_process_sct(r_master0_r_Pop_mioi_irdy_master_process_sct),
      .r_master0_r_Pop_mioi_ivld(r_master0_r_Pop_mioi_ivld)
    );
  scatter_gather_dma_master_process_r_master0_r_Pop_mioi_r_master0_r_Pop_mio_wait_dp
      scatter_gather_dma_master_process_r_master0_r_Pop_mioi_r_master0_r_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .r_master0_r_Pop_mioi_oswt_unreg(r_master0_r_Pop_mioi_oswt_unreg),
      .r_master0_r_Pop_mioi_bawt(r_master0_r_Pop_mioi_bawt),
      .r_master0_r_Pop_mioi_wen_comp(r_master0_r_Pop_mioi_wen_comp),
      .r_master0_r_Pop_mioi_idat_mxwt(r_master0_r_Pop_mioi_idat_mxwt_pconst),
      .r_master0_r_Pop_mioi_biwt(r_master0_r_Pop_mioi_biwt),
      .r_master0_r_Pop_mioi_bdwt(r_master0_r_Pop_mioi_bdwt),
      .r_master0_r_Pop_mioi_idat(r_master0_r_Pop_mioi_idat)
    );
  assign r_master0_r_Pop_mioi_idat_mxwt = r_master0_r_Pop_mioi_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi (
  clk, rst_bar, w_segment0_ex_aw_chan_vld, w_segment0_ex_aw_chan_rdy, w_segment0_ex_aw_chan_dat,
      master_process_wen, w_segment0_ex_aw_chan_Push_mioi_oswt, w_segment0_ex_aw_chan_Push_mioi_wen_comp,
      w_segment0_ex_aw_chan_Push_mioi_m_addr_rsc_dat_master_process, w_segment0_ex_aw_chan_Push_mioi_m_ex_len_rsc_dat_master_process,
      w_segment0_ex_aw_chan_Push_mioi_oswt_pff
);
  input clk;
  input rst_bar;
  output w_segment0_ex_aw_chan_vld;
  input w_segment0_ex_aw_chan_rdy;
  output [75:0] w_segment0_ex_aw_chan_dat;
  input master_process_wen;
  input w_segment0_ex_aw_chan_Push_mioi_oswt;
  output w_segment0_ex_aw_chan_Push_mioi_wen_comp;
  input [31:0] w_segment0_ex_aw_chan_Push_mioi_m_addr_rsc_dat_master_process;
  input [31:0] w_segment0_ex_aw_chan_Push_mioi_m_ex_len_rsc_dat_master_process;
  input w_segment0_ex_aw_chan_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire w_segment0_ex_aw_chan_Push_mioi_biwt;
  wire w_segment0_ex_aw_chan_Push_mioi_bdwt;
  wire w_segment0_ex_aw_chan_Push_mioi_bcwt;
  wire w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  wire w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_aw_payload_Connections_SYN_PORT_Push
      w_segment0_ex_aw_chan_Push_mioi (
      .this_vld(w_segment0_ex_aw_chan_vld),
      .this_rdy(w_segment0_ex_aw_chan_rdy),
      .this_dat(w_segment0_ex_aw_chan_dat),
      .m_addr_rsc_dat(w_segment0_ex_aw_chan_Push_mioi_m_addr_rsc_dat_master_process),
      .m_ex_len_rsc_dat(w_segment0_ex_aw_chan_Push_mioi_m_ex_len_rsc_dat_master_process),
      .ccs_ccore_start_rsc_dat(w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .ccs_ccore_done_sync_vld(w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_w_segment0_ex_aw_chan_Push_mio_wait_ctrl
      scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_w_segment0_ex_aw_chan_Push_mio_wait_ctrl_inst
      (
      .master_process_wen(master_process_wen),
      .w_segment0_ex_aw_chan_Push_mioi_oswt(w_segment0_ex_aw_chan_Push_mioi_oswt),
      .w_segment0_ex_aw_chan_Push_mioi_biwt(w_segment0_ex_aw_chan_Push_mioi_biwt),
      .w_segment0_ex_aw_chan_Push_mioi_bdwt(w_segment0_ex_aw_chan_Push_mioi_bdwt),
      .w_segment0_ex_aw_chan_Push_mioi_bcwt(w_segment0_ex_aw_chan_Push_mioi_bcwt),
      .w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct(w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_done_sync_vld(w_segment0_ex_aw_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .w_segment0_ex_aw_chan_Push_mioi_oswt_pff(w_segment0_ex_aw_chan_Push_mioi_oswt_pff)
    );
  scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_w_segment0_ex_aw_chan_Push_mio_wait_dp
      scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_w_segment0_ex_aw_chan_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_segment0_ex_aw_chan_Push_mioi_oswt(w_segment0_ex_aw_chan_Push_mioi_oswt),
      .w_segment0_ex_aw_chan_Push_mioi_wen_comp(w_segment0_ex_aw_chan_Push_mioi_wen_comp),
      .w_segment0_ex_aw_chan_Push_mioi_biwt(w_segment0_ex_aw_chan_Push_mioi_biwt),
      .w_segment0_ex_aw_chan_Push_mioi_bdwt(w_segment0_ex_aw_chan_Push_mioi_bdwt),
      .w_segment0_ex_aw_chan_Push_mioi_bcwt(w_segment0_ex_aw_chan_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi (
  clk, rst_bar, r_segment0_ex_ar_chan_vld, r_segment0_ex_ar_chan_rdy, r_segment0_ex_ar_chan_dat,
      master_process_wen, r_segment0_ex_ar_chan_Push_mioi_oswt, r_segment0_ex_ar_chan_Push_mioi_wen_comp,
      r_segment0_ex_ar_chan_Push_mioi_m_addr_rsc_dat_master_process, r_segment0_ex_ar_chan_Push_mioi_m_ex_len_rsc_dat_master_process,
      r_segment0_ex_ar_chan_Push_mioi_oswt_pff
);
  input clk;
  input rst_bar;
  output r_segment0_ex_ar_chan_vld;
  input r_segment0_ex_ar_chan_rdy;
  output [75:0] r_segment0_ex_ar_chan_dat;
  input master_process_wen;
  input r_segment0_ex_ar_chan_Push_mioi_oswt;
  output r_segment0_ex_ar_chan_Push_mioi_wen_comp;
  input [31:0] r_segment0_ex_ar_chan_Push_mioi_m_addr_rsc_dat_master_process;
  input [31:0] r_segment0_ex_ar_chan_Push_mioi_m_ex_len_rsc_dat_master_process;
  input r_segment0_ex_ar_chan_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire r_segment0_ex_ar_chan_Push_mioi_biwt;
  wire r_segment0_ex_ar_chan_Push_mioi_bdwt;
  wire r_segment0_ex_ar_chan_Push_mioi_bcwt;
  wire r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  wire r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_axi_axi4_segment_axi_cfg_standard_ex_ar_payload_Connections_SYN_PORT_Push
      r_segment0_ex_ar_chan_Push_mioi (
      .this_vld(r_segment0_ex_ar_chan_vld),
      .this_rdy(r_segment0_ex_ar_chan_rdy),
      .this_dat(r_segment0_ex_ar_chan_dat),
      .m_addr_rsc_dat(r_segment0_ex_ar_chan_Push_mioi_m_addr_rsc_dat_master_process),
      .m_ex_len_rsc_dat(r_segment0_ex_ar_chan_Push_mioi_m_ex_len_rsc_dat_master_process),
      .ccs_ccore_start_rsc_dat(r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .ccs_ccore_done_sync_vld(r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_r_segment0_ex_ar_chan_Push_mio_wait_ctrl
      scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_r_segment0_ex_ar_chan_Push_mio_wait_ctrl_inst
      (
      .master_process_wen(master_process_wen),
      .r_segment0_ex_ar_chan_Push_mioi_oswt(r_segment0_ex_ar_chan_Push_mioi_oswt),
      .r_segment0_ex_ar_chan_Push_mioi_biwt(r_segment0_ex_ar_chan_Push_mioi_biwt),
      .r_segment0_ex_ar_chan_Push_mioi_bdwt(r_segment0_ex_ar_chan_Push_mioi_bdwt),
      .r_segment0_ex_ar_chan_Push_mioi_bcwt(r_segment0_ex_ar_chan_Push_mioi_bcwt),
      .r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct(r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_done_sync_vld(r_segment0_ex_ar_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .r_segment0_ex_ar_chan_Push_mioi_oswt_pff(r_segment0_ex_ar_chan_Push_mioi_oswt_pff)
    );
  scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_r_segment0_ex_ar_chan_Push_mio_wait_dp
      scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_r_segment0_ex_ar_chan_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .r_segment0_ex_ar_chan_Push_mioi_oswt(r_segment0_ex_ar_chan_Push_mioi_oswt),
      .r_segment0_ex_ar_chan_Push_mioi_wen_comp(r_segment0_ex_ar_chan_Push_mioi_wen_comp),
      .r_segment0_ex_ar_chan_Push_mioi_biwt(r_segment0_ex_ar_chan_Push_mioi_biwt),
      .r_segment0_ex_ar_chan_Push_mioi_bdwt(r_segment0_ex_ar_chan_Push_mioi_bdwt),
      .r_segment0_ex_ar_chan_Push_mioi_bcwt(r_segment0_ex_ar_chan_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi (
  clk, rst_bar, dma_cmd_chan_vld, dma_cmd_chan_rdy, dma_cmd_chan_dat, master_process_wen,
      dma_cmd_chan_Pop_mioi_oswt, dma_cmd_chan_Pop_mioi_wen_comp, dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt,
      dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt, dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt,
      dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt, dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt,
      dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt, dma_cmd_chan_Pop_mioi_oswt_pff
);
  input clk;
  input rst_bar;
  input dma_cmd_chan_vld;
  output dma_cmd_chan_rdy;
  input [175:0] dma_cmd_chan_dat;
  input master_process_wen;
  input dma_cmd_chan_Pop_mioi_oswt;
  output dma_cmd_chan_Pop_mioi_wen_comp;
  output [31:0] dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt;
  output [31:0] dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt;
  output [31:0] dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt;
  output [31:0] dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt;
  output [15:0] dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt;
  output [15:0] dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt;
  input dma_cmd_chan_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire dma_cmd_chan_Pop_mioi_biwt;
  wire dma_cmd_chan_Pop_mioi_bdwt;
  wire dma_cmd_chan_Pop_mioi_bcwt;
  wire [31:0] dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z;
  wire [31:0] dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z;
  wire [31:0] dma_cmd_chan_Pop_mioi_return_total_len_rsc_z;
  wire [31:0] dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z;
  wire [15:0] dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z;
  wire [15:0] dma_cmd_chan_Pop_mioi_return_scatter_groups_rsc_z;
  wire [15:0] dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z;
  wire dma_cmd_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct;
  wire dma_cmd_chan_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_dma_cmd_Connections_SYN_PORT_Pop  dma_cmd_chan_Pop_mioi
      (
      .this_vld(dma_cmd_chan_vld),
      .this_rdy(dma_cmd_chan_rdy),
      .this_dat(dma_cmd_chan_dat),
      .return_ar_addr_rsc_z(dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z),
      .return_aw_addr_rsc_z(dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z),
      .return_total_len_rsc_z(dma_cmd_chan_Pop_mioi_return_total_len_rsc_z),
      .return_scatter_stride_rsc_z(dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z),
      .return_scatter_len_rsc_z(dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z),
      .return_scatter_groups_rsc_z(dma_cmd_chan_Pop_mioi_return_scatter_groups_rsc_z),
      .return_dma_mode_rsc_z(dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z),
      .ccs_ccore_start_rsc_dat(dma_cmd_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .ccs_ccore_done_sync_vld(dma_cmd_chan_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_dma_cmd_chan_Pop_mio_wait_ctrl
      scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_dma_cmd_chan_Pop_mio_wait_ctrl_inst
      (
      .master_process_wen(master_process_wen),
      .dma_cmd_chan_Pop_mioi_oswt(dma_cmd_chan_Pop_mioi_oswt),
      .dma_cmd_chan_Pop_mioi_biwt(dma_cmd_chan_Pop_mioi_biwt),
      .dma_cmd_chan_Pop_mioi_bdwt(dma_cmd_chan_Pop_mioi_bdwt),
      .dma_cmd_chan_Pop_mioi_bcwt(dma_cmd_chan_Pop_mioi_bcwt),
      .dma_cmd_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct(dma_cmd_chan_Pop_mioi_ccs_ccore_start_rsc_dat_master_process_sct),
      .dma_cmd_chan_Pop_mioi_ccs_ccore_done_sync_vld(dma_cmd_chan_Pop_mioi_ccs_ccore_done_sync_vld),
      .dma_cmd_chan_Pop_mioi_oswt_pff(dma_cmd_chan_Pop_mioi_oswt_pff)
    );
  scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_dma_cmd_chan_Pop_mio_wait_dp
      scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_dma_cmd_chan_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .dma_cmd_chan_Pop_mioi_oswt(dma_cmd_chan_Pop_mioi_oswt),
      .dma_cmd_chan_Pop_mioi_wen_comp(dma_cmd_chan_Pop_mioi_wen_comp),
      .dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_biwt(dma_cmd_chan_Pop_mioi_biwt),
      .dma_cmd_chan_Pop_mioi_bdwt(dma_cmd_chan_Pop_mioi_bdwt),
      .dma_cmd_chan_Pop_mioi_bcwt(dma_cmd_chan_Pop_mioi_bcwt),
      .dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z(dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z),
      .dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z(dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z),
      .dma_cmd_chan_Pop_mioi_return_total_len_rsc_z(dma_cmd_chan_Pop_mioi_return_total_len_rsc_z),
      .dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z(dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z),
      .dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z(dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z),
      .dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z(dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_w_slave0_b_Push_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_w_slave0_b_Push_mioi (
  clk, rst_bar, w_slave0_b_vld, w_slave0_b_rdy, w_slave0_b_dat, slave_process_wen,
      w_slave0_b_Push_mioi_oswt, w_slave0_b_Push_mioi_wen_comp, w_slave0_b_Push_mioi_idat_slave_process
);
  input clk;
  input rst_bar;
  output w_slave0_b_vld;
  input w_slave0_b_rdy;
  output [1:0] w_slave0_b_dat;
  input slave_process_wen;
  input w_slave0_b_Push_mioi_oswt;
  output w_slave0_b_Push_mioi_wen_comp;
  input [1:0] w_slave0_b_Push_mioi_idat_slave_process;


  // Interconnect Declarations
  wire w_slave0_b_Push_mioi_biwt;
  wire w_slave0_b_Push_mioi_bdwt;
  wire w_slave0_b_Push_mioi_bcwt;
  wire [1:0] w_slave0_b_Push_mioi_idat;
  wire w_slave0_b_Push_mioi_ivld_slave_process_sct;
  wire w_slave0_b_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  wire [1:0] nl_scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_dp_inst_w_slave0_b_Push_mioi_idat_slave_process;
  assign nl_scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_dp_inst_w_slave0_b_Push_mioi_idat_slave_process
      = {(w_slave0_b_Push_mioi_idat_slave_process[1]) , 1'b0};
  ccs_conn_out_wait_v1 #(.width(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) w_slave0_b_Push_mioi (
      .vld(w_slave0_b_vld),
      .rdy(w_slave0_b_rdy),
      .dat(w_slave0_b_dat),
      .idat(w_slave0_b_Push_mioi_idat),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1),
      .ivld(w_slave0_b_Push_mioi_ivld_slave_process_sct),
      .irdy(w_slave0_b_Push_mioi_irdy)
    );
  scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_ctrl
      scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_ctrl_inst
      (
      .slave_process_wen(slave_process_wen),
      .w_slave0_b_Push_mioi_oswt(w_slave0_b_Push_mioi_oswt),
      .w_slave0_b_Push_mioi_biwt(w_slave0_b_Push_mioi_biwt),
      .w_slave0_b_Push_mioi_bdwt(w_slave0_b_Push_mioi_bdwt),
      .w_slave0_b_Push_mioi_bcwt(w_slave0_b_Push_mioi_bcwt),
      .w_slave0_b_Push_mioi_ivld_slave_process_sct(w_slave0_b_Push_mioi_ivld_slave_process_sct),
      .w_slave0_b_Push_mioi_irdy(w_slave0_b_Push_mioi_irdy)
    );
  scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_dp
      scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_slave0_b_Push_mioi_oswt(w_slave0_b_Push_mioi_oswt),
      .w_slave0_b_Push_mioi_wen_comp(w_slave0_b_Push_mioi_wen_comp),
      .w_slave0_b_Push_mioi_idat_slave_process(nl_scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_w_slave0_b_Push_mio_wait_dp_inst_w_slave0_b_Push_mioi_idat_slave_process[1:0]),
      .w_slave0_b_Push_mioi_biwt(w_slave0_b_Push_mioi_biwt),
      .w_slave0_b_Push_mioi_bdwt(w_slave0_b_Push_mioi_bdwt),
      .w_slave0_b_Push_mioi_bcwt(w_slave0_b_Push_mioi_bcwt),
      .w_slave0_b_Push_mioi_idat(w_slave0_b_Push_mioi_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi (
  clk, rst_bar, dma_cmd_chan_vld, dma_cmd_chan_rdy, dma_cmd_chan_dat, slave_process_wen,
      dma_cmd_chan_Push_mioi_oswt, dma_cmd_chan_Push_mioi_wen_comp, dma_cmd_chan_Push_mioi_m_ar_addr_rsc_dat_slave_process,
      dma_cmd_chan_Push_mioi_m_aw_addr_rsc_dat_slave_process, dma_cmd_chan_Push_mioi_m_total_len_rsc_dat_slave_process,
      dma_cmd_chan_Push_mioi_m_scatter_stride_rsc_dat_slave_process, dma_cmd_chan_Push_mioi_m_scatter_len_rsc_dat_slave_process,
      dma_cmd_chan_Push_mioi_m_scatter_groups_rsc_dat_slave_process, dma_cmd_chan_Push_mioi_m_dma_mode_rsc_dat_slave_process,
      dma_cmd_chan_Push_mioi_oswt_pff
);
  input clk;
  input rst_bar;
  output dma_cmd_chan_vld;
  input dma_cmd_chan_rdy;
  output [175:0] dma_cmd_chan_dat;
  input slave_process_wen;
  input dma_cmd_chan_Push_mioi_oswt;
  output dma_cmd_chan_Push_mioi_wen_comp;
  input [31:0] dma_cmd_chan_Push_mioi_m_ar_addr_rsc_dat_slave_process;
  input [31:0] dma_cmd_chan_Push_mioi_m_aw_addr_rsc_dat_slave_process;
  input [31:0] dma_cmd_chan_Push_mioi_m_total_len_rsc_dat_slave_process;
  input [31:0] dma_cmd_chan_Push_mioi_m_scatter_stride_rsc_dat_slave_process;
  input [15:0] dma_cmd_chan_Push_mioi_m_scatter_len_rsc_dat_slave_process;
  input [15:0] dma_cmd_chan_Push_mioi_m_scatter_groups_rsc_dat_slave_process;
  input [15:0] dma_cmd_chan_Push_mioi_m_dma_mode_rsc_dat_slave_process;
  input dma_cmd_chan_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire dma_cmd_chan_Push_mioi_biwt;
  wire dma_cmd_chan_Push_mioi_bdwt;
  wire dma_cmd_chan_Push_mioi_bcwt;
  wire dma_cmd_chan_Push_mioi_ccs_ccore_start_rsc_dat_slave_process_sct;
  wire dma_cmd_chan_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_dma_cmd_Connections_SYN_PORT_Push  dma_cmd_chan_Push_mioi
      (
      .this_vld(dma_cmd_chan_vld),
      .this_rdy(dma_cmd_chan_rdy),
      .this_dat(dma_cmd_chan_dat),
      .m_ar_addr_rsc_dat(dma_cmd_chan_Push_mioi_m_ar_addr_rsc_dat_slave_process),
      .m_aw_addr_rsc_dat(dma_cmd_chan_Push_mioi_m_aw_addr_rsc_dat_slave_process),
      .m_total_len_rsc_dat(dma_cmd_chan_Push_mioi_m_total_len_rsc_dat_slave_process),
      .m_scatter_stride_rsc_dat(dma_cmd_chan_Push_mioi_m_scatter_stride_rsc_dat_slave_process),
      .m_scatter_len_rsc_dat(dma_cmd_chan_Push_mioi_m_scatter_len_rsc_dat_slave_process),
      .m_scatter_groups_rsc_dat(dma_cmd_chan_Push_mioi_m_scatter_groups_rsc_dat_slave_process),
      .m_dma_mode_rsc_dat(dma_cmd_chan_Push_mioi_m_dma_mode_rsc_dat_slave_process),
      .ccs_ccore_start_rsc_dat(dma_cmd_chan_Push_mioi_ccs_ccore_start_rsc_dat_slave_process_sct),
      .ccs_ccore_done_sync_vld(dma_cmd_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_dma_cmd_chan_Push_mio_wait_ctrl
      scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_dma_cmd_chan_Push_mio_wait_ctrl_inst
      (
      .slave_process_wen(slave_process_wen),
      .dma_cmd_chan_Push_mioi_oswt(dma_cmd_chan_Push_mioi_oswt),
      .dma_cmd_chan_Push_mioi_biwt(dma_cmd_chan_Push_mioi_biwt),
      .dma_cmd_chan_Push_mioi_bdwt(dma_cmd_chan_Push_mioi_bdwt),
      .dma_cmd_chan_Push_mioi_bcwt(dma_cmd_chan_Push_mioi_bcwt),
      .dma_cmd_chan_Push_mioi_ccs_ccore_start_rsc_dat_slave_process_sct(dma_cmd_chan_Push_mioi_ccs_ccore_start_rsc_dat_slave_process_sct),
      .dma_cmd_chan_Push_mioi_ccs_ccore_done_sync_vld(dma_cmd_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_cmd_chan_Push_mioi_oswt_pff(dma_cmd_chan_Push_mioi_oswt_pff)
    );
  scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_dma_cmd_chan_Push_mio_wait_dp
      scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_dma_cmd_chan_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .dma_cmd_chan_Push_mioi_oswt(dma_cmd_chan_Push_mioi_oswt),
      .dma_cmd_chan_Push_mioi_wen_comp(dma_cmd_chan_Push_mioi_wen_comp),
      .dma_cmd_chan_Push_mioi_biwt(dma_cmd_chan_Push_mioi_biwt),
      .dma_cmd_chan_Push_mioi_bdwt(dma_cmd_chan_Push_mioi_bdwt),
      .dma_cmd_chan_Push_mioi_bcwt(dma_cmd_chan_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi (
  clk, rst_bar, w_slave0_w_vld, w_slave0_w_rdy, w_slave0_w_dat, slave_process_wen,
      w_slave0_w_Pop_mioi_oswt, w_slave0_w_Pop_mioi_wen_comp, w_slave0_w_Pop_mioi_idat_mxwt
);
  input clk;
  input rst_bar;
  input w_slave0_w_vld;
  output w_slave0_w_rdy;
  input [31:0] w_slave0_w_dat;
  input slave_process_wen;
  input w_slave0_w_Pop_mioi_oswt;
  output w_slave0_w_Pop_mioi_wen_comp;
  output [31:0] w_slave0_w_Pop_mioi_idat_mxwt;


  // Interconnect Declarations
  wire w_slave0_w_Pop_mioi_biwt;
  wire w_slave0_w_Pop_mioi_bdwt;
  wire w_slave0_w_Pop_mioi_bcwt;
  wire [31:0] w_slave0_w_Pop_mioi_idat;
  wire w_slave0_w_Pop_mioi_irdy_slave_process_sct;
  wire w_slave0_w_Pop_mioi_ivld;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_in_wait_v1 #(.width(32'sd32),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) w_slave0_w_Pop_mioi (
      .vld(w_slave0_w_vld),
      .rdy(w_slave0_w_rdy),
      .dat(w_slave0_w_dat),
      .idat(w_slave0_w_Pop_mioi_idat),
      .irdy(w_slave0_w_Pop_mioi_irdy_slave_process_sct),
      .ivld(w_slave0_w_Pop_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1)
    );
  scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi_w_slave0_w_Pop_mio_wait_ctrl
      scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi_w_slave0_w_Pop_mio_wait_ctrl_inst
      (
      .slave_process_wen(slave_process_wen),
      .w_slave0_w_Pop_mioi_oswt(w_slave0_w_Pop_mioi_oswt),
      .w_slave0_w_Pop_mioi_biwt(w_slave0_w_Pop_mioi_biwt),
      .w_slave0_w_Pop_mioi_bdwt(w_slave0_w_Pop_mioi_bdwt),
      .w_slave0_w_Pop_mioi_bcwt(w_slave0_w_Pop_mioi_bcwt),
      .w_slave0_w_Pop_mioi_irdy_slave_process_sct(w_slave0_w_Pop_mioi_irdy_slave_process_sct),
      .w_slave0_w_Pop_mioi_ivld(w_slave0_w_Pop_mioi_ivld)
    );
  scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi_w_slave0_w_Pop_mio_wait_dp
      scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi_w_slave0_w_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_slave0_w_Pop_mioi_oswt(w_slave0_w_Pop_mioi_oswt),
      .w_slave0_w_Pop_mioi_wen_comp(w_slave0_w_Pop_mioi_wen_comp),
      .w_slave0_w_Pop_mioi_idat_mxwt(w_slave0_w_Pop_mioi_idat_mxwt),
      .w_slave0_w_Pop_mioi_biwt(w_slave0_w_Pop_mioi_biwt),
      .w_slave0_w_Pop_mioi_bdwt(w_slave0_w_Pop_mioi_bdwt),
      .w_slave0_w_Pop_mioi_bcwt(w_slave0_w_Pop_mioi_bcwt),
      .w_slave0_w_Pop_mioi_idat(w_slave0_w_Pop_mioi_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi (
  clk, rst_bar, w_slave0_aw_vld, w_slave0_aw_rdy, w_slave0_aw_dat, slave_process_wen,
      w_slave0_aw_Pop_mioi_oswt, w_slave0_aw_Pop_mioi_wen_comp, w_slave0_aw_Pop_mioi_idat_mxwt
);
  input clk;
  input rst_bar;
  input w_slave0_aw_vld;
  output w_slave0_aw_rdy;
  input [31:0] w_slave0_aw_dat;
  input slave_process_wen;
  input w_slave0_aw_Pop_mioi_oswt;
  output w_slave0_aw_Pop_mioi_wen_comp;
  output [31:0] w_slave0_aw_Pop_mioi_idat_mxwt;


  // Interconnect Declarations
  wire w_slave0_aw_Pop_mioi_biwt;
  wire w_slave0_aw_Pop_mioi_bdwt;
  wire w_slave0_aw_Pop_mioi_bcwt;
  wire [31:0] w_slave0_aw_Pop_mioi_idat;
  wire w_slave0_aw_Pop_mioi_irdy_slave_process_sct;
  wire w_slave0_aw_Pop_mioi_ivld;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_in_wait_v1 #(.width(32'sd32),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) w_slave0_aw_Pop_mioi (
      .vld(w_slave0_aw_vld),
      .rdy(w_slave0_aw_rdy),
      .dat(w_slave0_aw_dat),
      .idat(w_slave0_aw_Pop_mioi_idat),
      .irdy(w_slave0_aw_Pop_mioi_irdy_slave_process_sct),
      .ivld(w_slave0_aw_Pop_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1)
    );
  scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi_w_slave0_aw_Pop_mio_wait_ctrl
      scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi_w_slave0_aw_Pop_mio_wait_ctrl_inst
      (
      .slave_process_wen(slave_process_wen),
      .w_slave0_aw_Pop_mioi_oswt(w_slave0_aw_Pop_mioi_oswt),
      .w_slave0_aw_Pop_mioi_biwt(w_slave0_aw_Pop_mioi_biwt),
      .w_slave0_aw_Pop_mioi_bdwt(w_slave0_aw_Pop_mioi_bdwt),
      .w_slave0_aw_Pop_mioi_bcwt(w_slave0_aw_Pop_mioi_bcwt),
      .w_slave0_aw_Pop_mioi_irdy_slave_process_sct(w_slave0_aw_Pop_mioi_irdy_slave_process_sct),
      .w_slave0_aw_Pop_mioi_ivld(w_slave0_aw_Pop_mioi_ivld)
    );
  scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi_w_slave0_aw_Pop_mio_wait_dp
      scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi_w_slave0_aw_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_slave0_aw_Pop_mioi_oswt(w_slave0_aw_Pop_mioi_oswt),
      .w_slave0_aw_Pop_mioi_wen_comp(w_slave0_aw_Pop_mioi_wen_comp),
      .w_slave0_aw_Pop_mioi_idat_mxwt(w_slave0_aw_Pop_mioi_idat_mxwt),
      .w_slave0_aw_Pop_mioi_biwt(w_slave0_aw_Pop_mioi_biwt),
      .w_slave0_aw_Pop_mioi_bdwt(w_slave0_aw_Pop_mioi_bdwt),
      .w_slave0_aw_Pop_mioi_bcwt(w_slave0_aw_Pop_mioi_bcwt),
      .w_slave0_aw_Pop_mioi_idat(w_slave0_aw_Pop_mioi_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi (
  clk, rst_bar, b_chan_vld, b_chan_rdy, b_chan_dat, b_chan_Push_mioi_oswt_unreg,
      b_process_wen, b_process_wten, b_chan_Push_mioi_bawt, b_chan_Push_mioi_iswt0,
      b_chan_Push_mioi_wen_comp, b_chan_Push_mioi_idat
);
  input clk;
  input rst_bar;
  output b_chan_vld;
  input b_chan_rdy;
  output [5:0] b_chan_dat;
  input b_chan_Push_mioi_oswt_unreg;
  input b_process_wen;
  input b_process_wten;
  output b_chan_Push_mioi_bawt;
  input b_chan_Push_mioi_iswt0;
  output b_chan_Push_mioi_wen_comp;
  input [5:0] b_chan_Push_mioi_idat;


  // Interconnect Declarations
  wire b_chan_Push_mioi_biwt;
  wire b_chan_Push_mioi_bdwt;
  wire b_chan_Push_mioi_ivld_b_process_sct;
  wire b_chan_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_out_wait_v1 #(.width(32'sd6),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) b_chan_Push_mioi (
      .vld(b_chan_vld),
      .rdy(b_chan_rdy),
      .dat(b_chan_dat),
      .idat(b_chan_Push_mioi_idat),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1),
      .ivld(b_chan_Push_mioi_ivld_b_process_sct),
      .irdy(b_chan_Push_mioi_irdy)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_b_chan_Push_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_b_chan_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .b_chan_Push_mioi_oswt_unreg(b_chan_Push_mioi_oswt_unreg),
      .b_process_wen(b_process_wen),
      .b_process_wten(b_process_wten),
      .b_chan_Push_mioi_iswt0(b_chan_Push_mioi_iswt0),
      .b_chan_Push_mioi_biwt(b_chan_Push_mioi_biwt),
      .b_chan_Push_mioi_bdwt(b_chan_Push_mioi_bdwt),
      .b_chan_Push_mioi_ivld_b_process_sct(b_chan_Push_mioi_ivld_b_process_sct),
      .b_chan_Push_mioi_irdy(b_chan_Push_mioi_irdy)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_b_chan_Push_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_b_chan_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .b_chan_Push_mioi_oswt_unreg(b_chan_Push_mioi_oswt_unreg),
      .b_chan_Push_mioi_bawt(b_chan_Push_mioi_bawt),
      .b_chan_Push_mioi_wen_comp(b_chan_Push_mioi_wen_comp),
      .b_chan_Push_mioi_biwt(b_chan_Push_mioi_biwt),
      .b_chan_Push_mioi_bdwt(b_chan_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi
    (
  clk, rst_bar, last_burst_chan_vld, last_burst_chan_rdy, last_burst_chan_dat, last_burst_chan_Pop_mioi_oswt_unreg,
      b_process_wen, b_process_wten, last_burst_chan_Pop_mioi_bawt, last_burst_chan_Pop_mioi_iswt0,
      last_burst_chan_Pop_mioi_wen_comp, last_burst_chan_Pop_mioi_return_rsc_z_mxwt,
      last_burst_chan_Pop_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  input last_burst_chan_vld;
  output last_burst_chan_rdy;
  input last_burst_chan_dat;
  input last_burst_chan_Pop_mioi_oswt_unreg;
  input b_process_wen;
  input b_process_wten;
  output last_burst_chan_Pop_mioi_bawt;
  input last_burst_chan_Pop_mioi_iswt0;
  output last_burst_chan_Pop_mioi_wen_comp;
  output last_burst_chan_Pop_mioi_return_rsc_z_mxwt;
  input last_burst_chan_Pop_mioi_iswt0_pff;


  // Interconnect Declarations
  wire last_burst_chan_Pop_mioi_biwt;
  wire last_burst_chan_Pop_mioi_bdwt;
  wire last_burst_chan_Pop_mioi_return_rsc_z;
  wire last_burst_chan_Pop_mioi_ccs_ccore_start_rsc_dat_b_process_sct;
  wire last_burst_chan_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_bool_Connections_SYN_PORT_Pop  last_burst_chan_Pop_mioi
      (
      .this_vld(last_burst_chan_vld),
      .this_rdy(last_burst_chan_rdy),
      .this_dat(last_burst_chan_dat),
      .return_rsc_z(last_burst_chan_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(last_burst_chan_Pop_mioi_ccs_ccore_start_rsc_dat_b_process_sct),
      .ccs_ccore_done_sync_vld(last_burst_chan_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi_last_burst_chan_Pop_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi_last_burst_chan_Pop_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_burst_chan_Pop_mioi_oswt_unreg(last_burst_chan_Pop_mioi_oswt_unreg),
      .b_process_wen(b_process_wen),
      .b_process_wten(b_process_wten),
      .last_burst_chan_Pop_mioi_iswt0(last_burst_chan_Pop_mioi_iswt0),
      .last_burst_chan_Pop_mioi_biwt(last_burst_chan_Pop_mioi_biwt),
      .last_burst_chan_Pop_mioi_bdwt(last_burst_chan_Pop_mioi_bdwt),
      .last_burst_chan_Pop_mioi_ccs_ccore_start_rsc_dat_b_process_sct(last_burst_chan_Pop_mioi_ccs_ccore_start_rsc_dat_b_process_sct),
      .last_burst_chan_Pop_mioi_ccs_ccore_done_sync_vld(last_burst_chan_Pop_mioi_ccs_ccore_done_sync_vld),
      .last_burst_chan_Pop_mioi_iswt0_pff(last_burst_chan_Pop_mioi_iswt0_pff)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi_last_burst_chan_Pop_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi_last_burst_chan_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_burst_chan_Pop_mioi_oswt_unreg(last_burst_chan_Pop_mioi_oswt_unreg),
      .last_burst_chan_Pop_mioi_bawt(last_burst_chan_Pop_mioi_bawt),
      .last_burst_chan_Pop_mioi_wen_comp(last_burst_chan_Pop_mioi_wen_comp),
      .last_burst_chan_Pop_mioi_return_rsc_z_mxwt(last_burst_chan_Pop_mioi_return_rsc_z_mxwt),
      .last_burst_chan_Pop_mioi_biwt(last_burst_chan_Pop_mioi_biwt),
      .last_burst_chan_Pop_mioi_bdwt(last_burst_chan_Pop_mioi_bdwt),
      .last_burst_chan_Pop_mioi_return_rsc_z(last_burst_chan_Pop_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi (
  clk, rst_bar, b_in_vld, b_in_rdy, b_in_dat, b_in_Pop_mioi_oswt_unreg, b_process_wen,
      b_process_wten, b_in_Pop_mioi_bawt, b_in_Pop_mioi_iswt0, b_in_Pop_mioi_wen_comp,
      b_in_Pop_mioi_idat_mxwt
);
  input clk;
  input rst_bar;
  input b_in_vld;
  output b_in_rdy;
  input [5:0] b_in_dat;
  input b_in_Pop_mioi_oswt_unreg;
  input b_process_wen;
  input b_process_wten;
  output b_in_Pop_mioi_bawt;
  input b_in_Pop_mioi_iswt0;
  output b_in_Pop_mioi_wen_comp;
  output [5:0] b_in_Pop_mioi_idat_mxwt;


  // Interconnect Declarations
  wire b_in_Pop_mioi_biwt;
  wire b_in_Pop_mioi_bdwt;
  wire [5:0] b_in_Pop_mioi_idat;
  wire b_in_Pop_mioi_irdy_b_process_sct;
  wire b_in_Pop_mioi_ivld;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_in_wait_v1 #(.width(32'sd6),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) b_in_Pop_mioi (
      .vld(b_in_vld),
      .rdy(b_in_rdy),
      .dat(b_in_dat),
      .idat(b_in_Pop_mioi_idat),
      .irdy(b_in_Pop_mioi_irdy_b_process_sct),
      .ivld(b_in_Pop_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi_b_in_Pop_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi_b_in_Pop_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .b_in_Pop_mioi_oswt_unreg(b_in_Pop_mioi_oswt_unreg),
      .b_process_wen(b_process_wen),
      .b_process_wten(b_process_wten),
      .b_in_Pop_mioi_iswt0(b_in_Pop_mioi_iswt0),
      .b_in_Pop_mioi_biwt(b_in_Pop_mioi_biwt),
      .b_in_Pop_mioi_bdwt(b_in_Pop_mioi_bdwt),
      .b_in_Pop_mioi_irdy_b_process_sct(b_in_Pop_mioi_irdy_b_process_sct),
      .b_in_Pop_mioi_ivld(b_in_Pop_mioi_ivld)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi_b_in_Pop_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi_b_in_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .b_in_Pop_mioi_oswt_unreg(b_in_Pop_mioi_oswt_unreg),
      .b_in_Pop_mioi_bawt(b_in_Pop_mioi_bawt),
      .b_in_Pop_mioi_wen_comp(b_in_Pop_mioi_wen_comp),
      .b_in_Pop_mioi_idat_mxwt(b_in_Pop_mioi_idat_mxwt),
      .b_in_Pop_mioi_biwt(b_in_Pop_mioi_biwt),
      .b_in_Pop_mioi_bdwt(b_in_Pop_mioi_bdwt),
      .b_in_Pop_mioi_idat(b_in_Pop_mioi_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi (
  clk, rst_bar, w_out_vld, w_out_rdy, w_out_dat, w_out_Push_mioi_oswt_unreg, w_process_wen,
      w_process_wten, w_out_Push_mioi_bawt, w_out_Push_mioi_iswt0, w_out_Push_mioi_wen_comp,
      w_out_Push_mioi_idat
);
  input clk;
  input rst_bar;
  output w_out_vld;
  input w_out_rdy;
  output [72:0] w_out_dat;
  input w_out_Push_mioi_oswt_unreg;
  input w_process_wen;
  input w_process_wten;
  output w_out_Push_mioi_bawt;
  input w_out_Push_mioi_iswt0;
  output w_out_Push_mioi_wen_comp;
  input [72:0] w_out_Push_mioi_idat;


  // Interconnect Declarations
  wire w_out_Push_mioi_biwt;
  wire w_out_Push_mioi_bdwt;
  wire w_out_Push_mioi_ivld_w_process_sct;
  wire w_out_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_out_wait_v1 #(.width(32'sd73),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) w_out_Push_mioi (
      .vld(w_out_vld),
      .rdy(w_out_rdy),
      .dat(w_out_dat),
      .idat(w_out_Push_mioi_idat),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1),
      .ivld(w_out_Push_mioi_ivld_w_process_sct),
      .irdy(w_out_Push_mioi_irdy)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_w_out_Push_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_w_out_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_out_Push_mioi_oswt_unreg(w_out_Push_mioi_oswt_unreg),
      .w_process_wen(w_process_wen),
      .w_process_wten(w_process_wten),
      .w_out_Push_mioi_iswt0(w_out_Push_mioi_iswt0),
      .w_out_Push_mioi_biwt(w_out_Push_mioi_biwt),
      .w_out_Push_mioi_bdwt(w_out_Push_mioi_bdwt),
      .w_out_Push_mioi_ivld_w_process_sct(w_out_Push_mioi_ivld_w_process_sct),
      .w_out_Push_mioi_irdy(w_out_Push_mioi_irdy)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_w_out_Push_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_w_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_out_Push_mioi_oswt_unreg(w_out_Push_mioi_oswt_unreg),
      .w_out_Push_mioi_bawt(w_out_Push_mioi_bawt),
      .w_out_Push_mioi_wen_comp(w_out_Push_mioi_wen_comp),
      .w_out_Push_mioi_biwt(w_out_Push_mioi_biwt),
      .w_out_Push_mioi_bdwt(w_out_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi
    (
  clk, rst_bar, last_bit_chan_vld, last_bit_chan_rdy, last_bit_chan_dat, last_bit_chan_Pop_mioi_oswt_unreg,
      w_process_wen, w_process_wten, last_bit_chan_Pop_mioi_bawt, last_bit_chan_Pop_mioi_iswt0,
      last_bit_chan_Pop_mioi_wen_comp, last_bit_chan_Pop_mioi_return_rsc_z_mxwt,
      last_bit_chan_Pop_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  input last_bit_chan_vld;
  output last_bit_chan_rdy;
  input last_bit_chan_dat;
  input last_bit_chan_Pop_mioi_oswt_unreg;
  input w_process_wen;
  input w_process_wten;
  output last_bit_chan_Pop_mioi_bawt;
  input last_bit_chan_Pop_mioi_iswt0;
  output last_bit_chan_Pop_mioi_wen_comp;
  output last_bit_chan_Pop_mioi_return_rsc_z_mxwt;
  input last_bit_chan_Pop_mioi_iswt0_pff;


  // Interconnect Declarations
  wire last_bit_chan_Pop_mioi_biwt;
  wire last_bit_chan_Pop_mioi_bdwt;
  wire last_bit_chan_Pop_mioi_return_rsc_z;
  wire last_bit_chan_Pop_mioi_ccs_ccore_start_rsc_dat_w_process_sct;
  wire last_bit_chan_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_bool_Connections_SYN_PORT_Pop  last_bit_chan_Pop_mioi
      (
      .this_vld(last_bit_chan_vld),
      .this_rdy(last_bit_chan_rdy),
      .this_dat(last_bit_chan_dat),
      .return_rsc_z(last_bit_chan_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(last_bit_chan_Pop_mioi_ccs_ccore_start_rsc_dat_w_process_sct),
      .ccs_ccore_done_sync_vld(last_bit_chan_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi_last_bit_chan_Pop_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi_last_bit_chan_Pop_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_bit_chan_Pop_mioi_oswt_unreg(last_bit_chan_Pop_mioi_oswt_unreg),
      .w_process_wen(w_process_wen),
      .w_process_wten(w_process_wten),
      .last_bit_chan_Pop_mioi_iswt0(last_bit_chan_Pop_mioi_iswt0),
      .last_bit_chan_Pop_mioi_biwt(last_bit_chan_Pop_mioi_biwt),
      .last_bit_chan_Pop_mioi_bdwt(last_bit_chan_Pop_mioi_bdwt),
      .last_bit_chan_Pop_mioi_ccs_ccore_start_rsc_dat_w_process_sct(last_bit_chan_Pop_mioi_ccs_ccore_start_rsc_dat_w_process_sct),
      .last_bit_chan_Pop_mioi_ccs_ccore_done_sync_vld(last_bit_chan_Pop_mioi_ccs_ccore_done_sync_vld),
      .last_bit_chan_Pop_mioi_iswt0_pff(last_bit_chan_Pop_mioi_iswt0_pff)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi_last_bit_chan_Pop_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi_last_bit_chan_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_bit_chan_Pop_mioi_oswt_unreg(last_bit_chan_Pop_mioi_oswt_unreg),
      .last_bit_chan_Pop_mioi_bawt(last_bit_chan_Pop_mioi_bawt),
      .last_bit_chan_Pop_mioi_wen_comp(last_bit_chan_Pop_mioi_wen_comp),
      .last_bit_chan_Pop_mioi_return_rsc_z_mxwt(last_bit_chan_Pop_mioi_return_rsc_z_mxwt),
      .last_bit_chan_Pop_mioi_biwt(last_bit_chan_Pop_mioi_biwt),
      .last_bit_chan_Pop_mioi_bdwt(last_bit_chan_Pop_mioi_bdwt),
      .last_bit_chan_Pop_mioi_return_rsc_z(last_bit_chan_Pop_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi (
  clk, rst_bar, w_chan_vld, w_chan_rdy, w_chan_dat, w_chan_Pop_mioi_oswt_unreg, w_process_wen,
      w_process_wten, w_chan_Pop_mioi_bawt, w_chan_Pop_mioi_iswt0, w_chan_Pop_mioi_wen_comp,
      w_chan_Pop_mioi_idat_mxwt
);
  input clk;
  input rst_bar;
  input w_chan_vld;
  output w_chan_rdy;
  input [72:0] w_chan_dat;
  input w_chan_Pop_mioi_oswt_unreg;
  input w_process_wen;
  input w_process_wten;
  output w_chan_Pop_mioi_bawt;
  input w_chan_Pop_mioi_iswt0;
  output w_chan_Pop_mioi_wen_comp;
  output [71:0] w_chan_Pop_mioi_idat_mxwt;


  // Interconnect Declarations
  wire w_chan_Pop_mioi_biwt;
  wire w_chan_Pop_mioi_bdwt;
  wire [72:0] w_chan_Pop_mioi_idat;
  wire w_chan_Pop_mioi_irdy_w_process_sct;
  wire w_chan_Pop_mioi_ivld;
  wire [71:0] w_chan_Pop_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_in_wait_v1 #(.width(32'sd73),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) w_chan_Pop_mioi (
      .vld(w_chan_vld),
      .rdy(w_chan_rdy),
      .dat(w_chan_dat),
      .idat(w_chan_Pop_mioi_idat),
      .irdy(w_chan_Pop_mioi_irdy_w_process_sct),
      .ivld(w_chan_Pop_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi_w_chan_Pop_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi_w_chan_Pop_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_chan_Pop_mioi_oswt_unreg(w_chan_Pop_mioi_oswt_unreg),
      .w_process_wen(w_process_wen),
      .w_process_wten(w_process_wten),
      .w_chan_Pop_mioi_iswt0(w_chan_Pop_mioi_iswt0),
      .w_chan_Pop_mioi_biwt(w_chan_Pop_mioi_biwt),
      .w_chan_Pop_mioi_bdwt(w_chan_Pop_mioi_bdwt),
      .w_chan_Pop_mioi_irdy_w_process_sct(w_chan_Pop_mioi_irdy_w_process_sct),
      .w_chan_Pop_mioi_ivld(w_chan_Pop_mioi_ivld)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi_w_chan_Pop_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi_w_chan_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_chan_Pop_mioi_oswt_unreg(w_chan_Pop_mioi_oswt_unreg),
      .w_chan_Pop_mioi_bawt(w_chan_Pop_mioi_bawt),
      .w_chan_Pop_mioi_wen_comp(w_chan_Pop_mioi_wen_comp),
      .w_chan_Pop_mioi_idat_mxwt(w_chan_Pop_mioi_idat_mxwt_pconst),
      .w_chan_Pop_mioi_biwt(w_chan_Pop_mioi_biwt),
      .w_chan_Pop_mioi_bdwt(w_chan_Pop_mioi_bdwt),
      .w_chan_Pop_mioi_idat(w_chan_Pop_mioi_idat)
    );
  assign w_chan_Pop_mioi_idat_mxwt = w_chan_Pop_mioi_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi
    (
  clk, rst_bar, last_burst_chan_vld, last_burst_chan_rdy, last_burst_chan_dat, ex_aw_process_wen,
      ex_aw_process_wten, last_burst_chan_Push_mioi_oswt_unreg, last_burst_chan_Push_mioi_bawt,
      last_burst_chan_Push_mioi_iswt0, last_burst_chan_Push_mioi_wen_comp, last_burst_chan_Push_mioi_m_rsc_dat,
      last_burst_chan_Push_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  output last_burst_chan_vld;
  input last_burst_chan_rdy;
  output last_burst_chan_dat;
  input ex_aw_process_wen;
  input ex_aw_process_wten;
  input last_burst_chan_Push_mioi_oswt_unreg;
  output last_burst_chan_Push_mioi_bawt;
  input last_burst_chan_Push_mioi_iswt0;
  output last_burst_chan_Push_mioi_wen_comp;
  input last_burst_chan_Push_mioi_m_rsc_dat;
  input last_burst_chan_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire last_burst_chan_Push_mioi_biwt;
  wire last_burst_chan_Push_mioi_bdwt;
  wire last_burst_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct;
  wire last_burst_chan_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_bool_Connections_SYN_PORT_Push  last_burst_chan_Push_mioi
      (
      .this_vld(last_burst_chan_vld),
      .this_rdy(last_burst_chan_rdy),
      .this_dat(last_burst_chan_dat),
      .m_rsc_dat(last_burst_chan_Push_mioi_m_rsc_dat),
      .ccs_ccore_start_rsc_dat(last_burst_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct),
      .ccs_ccore_done_sync_vld(last_burst_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_last_burst_chan_Push_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_last_burst_chan_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_aw_process_wen(ex_aw_process_wen),
      .ex_aw_process_wten(ex_aw_process_wten),
      .last_burst_chan_Push_mioi_oswt_unreg(last_burst_chan_Push_mioi_oswt_unreg),
      .last_burst_chan_Push_mioi_iswt0(last_burst_chan_Push_mioi_iswt0),
      .last_burst_chan_Push_mioi_biwt(last_burst_chan_Push_mioi_biwt),
      .last_burst_chan_Push_mioi_bdwt(last_burst_chan_Push_mioi_bdwt),
      .last_burst_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct(last_burst_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct),
      .last_burst_chan_Push_mioi_ccs_ccore_done_sync_vld(last_burst_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .last_burst_chan_Push_mioi_iswt0_pff(last_burst_chan_Push_mioi_iswt0_pff)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_last_burst_chan_Push_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_last_burst_chan_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_burst_chan_Push_mioi_oswt_unreg(last_burst_chan_Push_mioi_oswt_unreg),
      .last_burst_chan_Push_mioi_bawt(last_burst_chan_Push_mioi_bawt),
      .last_burst_chan_Push_mioi_wen_comp(last_burst_chan_Push_mioi_wen_comp),
      .last_burst_chan_Push_mioi_biwt(last_burst_chan_Push_mioi_biwt),
      .last_burst_chan_Push_mioi_bdwt(last_burst_chan_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi
    (
  clk, rst_bar, last_bit_chan_vld, last_bit_chan_rdy, last_bit_chan_dat, ex_aw_process_wen,
      ex_aw_process_wten, last_bit_chan_Push_mioi_oswt_unreg, last_bit_chan_Push_mioi_bawt,
      last_bit_chan_Push_mioi_iswt0, last_bit_chan_Push_mioi_wen_comp, last_bit_chan_Push_mioi_m_rsc_dat,
      last_bit_chan_Push_mioi_iswt0_pff
);
  input clk;
  input rst_bar;
  output last_bit_chan_vld;
  input last_bit_chan_rdy;
  output last_bit_chan_dat;
  input ex_aw_process_wen;
  input ex_aw_process_wten;
  input last_bit_chan_Push_mioi_oswt_unreg;
  output last_bit_chan_Push_mioi_bawt;
  input last_bit_chan_Push_mioi_iswt0;
  output last_bit_chan_Push_mioi_wen_comp;
  input last_bit_chan_Push_mioi_m_rsc_dat;
  input last_bit_chan_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire last_bit_chan_Push_mioi_biwt;
  wire last_bit_chan_Push_mioi_bdwt;
  wire last_bit_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct;
  wire last_bit_chan_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_bool_Connections_SYN_PORT_Push  last_bit_chan_Push_mioi
      (
      .this_vld(last_bit_chan_vld),
      .this_rdy(last_bit_chan_rdy),
      .this_dat(last_bit_chan_dat),
      .m_rsc_dat(last_bit_chan_Push_mioi_m_rsc_dat),
      .ccs_ccore_start_rsc_dat(last_bit_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct),
      .ccs_ccore_done_sync_vld(last_bit_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst_bar)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_last_bit_chan_Push_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_last_bit_chan_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_aw_process_wen(ex_aw_process_wen),
      .ex_aw_process_wten(ex_aw_process_wten),
      .last_bit_chan_Push_mioi_oswt_unreg(last_bit_chan_Push_mioi_oswt_unreg),
      .last_bit_chan_Push_mioi_iswt0(last_bit_chan_Push_mioi_iswt0),
      .last_bit_chan_Push_mioi_biwt(last_bit_chan_Push_mioi_biwt),
      .last_bit_chan_Push_mioi_bdwt(last_bit_chan_Push_mioi_bdwt),
      .last_bit_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct(last_bit_chan_Push_mioi_ccs_ccore_start_rsc_dat_ex_aw_process_sct),
      .last_bit_chan_Push_mioi_ccs_ccore_done_sync_vld(last_bit_chan_Push_mioi_ccs_ccore_done_sync_vld),
      .last_bit_chan_Push_mioi_iswt0_pff(last_bit_chan_Push_mioi_iswt0_pff)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_last_bit_chan_Push_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_last_bit_chan_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_bit_chan_Push_mioi_oswt_unreg(last_bit_chan_Push_mioi_oswt_unreg),
      .last_bit_chan_Push_mioi_bawt(last_bit_chan_Push_mioi_bawt),
      .last_bit_chan_Push_mioi_wen_comp(last_bit_chan_Push_mioi_wen_comp),
      .last_bit_chan_Push_mioi_biwt(last_bit_chan_Push_mioi_biwt),
      .last_bit_chan_Push_mioi_bdwt(last_bit_chan_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi
    (
  clk, rst_bar, aw_out_vld, aw_out_rdy, aw_out_dat, ex_aw_process_wen, ex_aw_process_wten,
      aw_out_Push_mioi_oswt_unreg, aw_out_Push_mioi_bawt, aw_out_Push_mioi_iswt0,
      aw_out_Push_mioi_wen_comp, aw_out_Push_mioi_idat
);
  input clk;
  input rst_bar;
  output aw_out_vld;
  input aw_out_rdy;
  output [43:0] aw_out_dat;
  input ex_aw_process_wen;
  input ex_aw_process_wten;
  input aw_out_Push_mioi_oswt_unreg;
  output aw_out_Push_mioi_bawt;
  input aw_out_Push_mioi_iswt0;
  output aw_out_Push_mioi_wen_comp;
  input [43:0] aw_out_Push_mioi_idat;


  // Interconnect Declarations
  wire aw_out_Push_mioi_biwt;
  wire aw_out_Push_mioi_bdwt;
  wire aw_out_Push_mioi_ivld_ex_aw_process_sct;
  wire aw_out_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_out_wait_v1 #(.width(32'sd44),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) aw_out_Push_mioi (
      .vld(aw_out_vld),
      .rdy(aw_out_rdy),
      .dat(aw_out_dat),
      .idat(aw_out_Push_mioi_idat),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1),
      .ivld(aw_out_Push_mioi_ivld_ex_aw_process_sct),
      .irdy(aw_out_Push_mioi_irdy)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_aw_out_Push_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_aw_out_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_aw_process_wen(ex_aw_process_wen),
      .ex_aw_process_wten(ex_aw_process_wten),
      .aw_out_Push_mioi_oswt_unreg(aw_out_Push_mioi_oswt_unreg),
      .aw_out_Push_mioi_iswt0(aw_out_Push_mioi_iswt0),
      .aw_out_Push_mioi_biwt(aw_out_Push_mioi_biwt),
      .aw_out_Push_mioi_bdwt(aw_out_Push_mioi_bdwt),
      .aw_out_Push_mioi_ivld_ex_aw_process_sct(aw_out_Push_mioi_ivld_ex_aw_process_sct),
      .aw_out_Push_mioi_irdy(aw_out_Push_mioi_irdy)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_aw_out_Push_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_aw_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .aw_out_Push_mioi_oswt_unreg(aw_out_Push_mioi_oswt_unreg),
      .aw_out_Push_mioi_bawt(aw_out_Push_mioi_bawt),
      .aw_out_Push_mioi_wen_comp(aw_out_Push_mioi_wen_comp),
      .aw_out_Push_mioi_biwt(aw_out_Push_mioi_biwt),
      .aw_out_Push_mioi_bdwt(aw_out_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi
    (
  clk, rst_bar, ex_aw_chan_vld, ex_aw_chan_rdy, ex_aw_chan_dat, ex_aw_process_wen,
      ex_aw_process_wten, ex_aw_chan_Pop_mioi_oswt_unreg, ex_aw_chan_Pop_mioi_bawt,
      ex_aw_chan_Pop_mioi_iswt0, ex_aw_chan_Pop_mioi_wen_comp, ex_aw_chan_Pop_mioi_idat_mxwt
);
  input clk;
  input rst_bar;
  input ex_aw_chan_vld;
  output ex_aw_chan_rdy;
  input [75:0] ex_aw_chan_dat;
  input ex_aw_process_wen;
  input ex_aw_process_wten;
  input ex_aw_chan_Pop_mioi_oswt_unreg;
  output ex_aw_chan_Pop_mioi_bawt;
  input ex_aw_chan_Pop_mioi_iswt0;
  output ex_aw_chan_Pop_mioi_wen_comp;
  output [67:0] ex_aw_chan_Pop_mioi_idat_mxwt;


  // Interconnect Declarations
  wire ex_aw_chan_Pop_mioi_biwt;
  wire ex_aw_chan_Pop_mioi_bdwt;
  wire [75:0] ex_aw_chan_Pop_mioi_idat;
  wire ex_aw_chan_Pop_mioi_irdy_ex_aw_process_sct;
  wire ex_aw_chan_Pop_mioi_ivld;
  wire [67:0] ex_aw_chan_Pop_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_in_wait_v1 #(.width(32'sd76),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ex_aw_chan_Pop_mioi (
      .vld(ex_aw_chan_vld),
      .rdy(ex_aw_chan_rdy),
      .dat(ex_aw_chan_dat),
      .idat(ex_aw_chan_Pop_mioi_idat),
      .irdy(ex_aw_chan_Pop_mioi_irdy_ex_aw_process_sct),
      .ivld(ex_aw_chan_Pop_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_ex_aw_chan_Pop_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_ex_aw_chan_Pop_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_aw_process_wen(ex_aw_process_wen),
      .ex_aw_process_wten(ex_aw_process_wten),
      .ex_aw_chan_Pop_mioi_oswt_unreg(ex_aw_chan_Pop_mioi_oswt_unreg),
      .ex_aw_chan_Pop_mioi_iswt0(ex_aw_chan_Pop_mioi_iswt0),
      .ex_aw_chan_Pop_mioi_biwt(ex_aw_chan_Pop_mioi_biwt),
      .ex_aw_chan_Pop_mioi_bdwt(ex_aw_chan_Pop_mioi_bdwt),
      .ex_aw_chan_Pop_mioi_irdy_ex_aw_process_sct(ex_aw_chan_Pop_mioi_irdy_ex_aw_process_sct),
      .ex_aw_chan_Pop_mioi_ivld(ex_aw_chan_Pop_mioi_ivld)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_ex_aw_chan_Pop_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_ex_aw_chan_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_aw_chan_Pop_mioi_oswt_unreg(ex_aw_chan_Pop_mioi_oswt_unreg),
      .ex_aw_chan_Pop_mioi_bawt(ex_aw_chan_Pop_mioi_bawt),
      .ex_aw_chan_Pop_mioi_wen_comp(ex_aw_chan_Pop_mioi_wen_comp),
      .ex_aw_chan_Pop_mioi_idat_mxwt(ex_aw_chan_Pop_mioi_idat_mxwt_pconst),
      .ex_aw_chan_Pop_mioi_biwt(ex_aw_chan_Pop_mioi_biwt),
      .ex_aw_chan_Pop_mioi_bdwt(ex_aw_chan_Pop_mioi_bdwt),
      .ex_aw_chan_Pop_mioi_idat(ex_aw_chan_Pop_mioi_idat)
    );
  assign ex_aw_chan_Pop_mioi_idat_mxwt = ex_aw_chan_Pop_mioi_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi
    (
  clk, rst_bar, ar_out_vld, ar_out_rdy, ar_out_dat, ex_ar_process_wen, ex_ar_process_wten,
      ar_out_Push_mioi_oswt_unreg, ar_out_Push_mioi_bawt, ar_out_Push_mioi_iswt0,
      ar_out_Push_mioi_wen_comp, ar_out_Push_mioi_idat
);
  input clk;
  input rst_bar;
  output ar_out_vld;
  input ar_out_rdy;
  output [43:0] ar_out_dat;
  input ex_ar_process_wen;
  input ex_ar_process_wten;
  input ar_out_Push_mioi_oswt_unreg;
  output ar_out_Push_mioi_bawt;
  input ar_out_Push_mioi_iswt0;
  output ar_out_Push_mioi_wen_comp;
  input [43:0] ar_out_Push_mioi_idat;


  // Interconnect Declarations
  wire ar_out_Push_mioi_biwt;
  wire ar_out_Push_mioi_bdwt;
  wire ar_out_Push_mioi_ivld_ex_ar_process_sct;
  wire ar_out_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_out_wait_v1 #(.width(32'sd44),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ar_out_Push_mioi (
      .vld(ar_out_vld),
      .rdy(ar_out_rdy),
      .dat(ar_out_dat),
      .idat(ar_out_Push_mioi_idat),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1),
      .ivld(ar_out_Push_mioi_ivld_ex_ar_process_sct),
      .irdy(ar_out_Push_mioi_irdy)
    );
  axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_ar_out_Push_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_ar_out_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_ar_process_wen(ex_ar_process_wen),
      .ex_ar_process_wten(ex_ar_process_wten),
      .ar_out_Push_mioi_oswt_unreg(ar_out_Push_mioi_oswt_unreg),
      .ar_out_Push_mioi_iswt0(ar_out_Push_mioi_iswt0),
      .ar_out_Push_mioi_biwt(ar_out_Push_mioi_biwt),
      .ar_out_Push_mioi_bdwt(ar_out_Push_mioi_bdwt),
      .ar_out_Push_mioi_ivld_ex_ar_process_sct(ar_out_Push_mioi_ivld_ex_ar_process_sct),
      .ar_out_Push_mioi_irdy(ar_out_Push_mioi_irdy)
    );
  axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_ar_out_Push_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_ar_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ar_out_Push_mioi_oswt_unreg(ar_out_Push_mioi_oswt_unreg),
      .ar_out_Push_mioi_bawt(ar_out_Push_mioi_bawt),
      .ar_out_Push_mioi_wen_comp(ar_out_Push_mioi_wen_comp),
      .ar_out_Push_mioi_biwt(ar_out_Push_mioi_biwt),
      .ar_out_Push_mioi_bdwt(ar_out_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi
    (
  clk, rst_bar, ex_ar_chan_vld, ex_ar_chan_rdy, ex_ar_chan_dat, ex_ar_process_wen,
      ex_ar_process_wten, ex_ar_chan_Pop_mioi_oswt_unreg, ex_ar_chan_Pop_mioi_bawt,
      ex_ar_chan_Pop_mioi_iswt0, ex_ar_chan_Pop_mioi_wen_comp, ex_ar_chan_Pop_mioi_idat_mxwt
);
  input clk;
  input rst_bar;
  input ex_ar_chan_vld;
  output ex_ar_chan_rdy;
  input [75:0] ex_ar_chan_dat;
  input ex_ar_process_wen;
  input ex_ar_process_wten;
  input ex_ar_chan_Pop_mioi_oswt_unreg;
  output ex_ar_chan_Pop_mioi_bawt;
  input ex_ar_chan_Pop_mioi_iswt0;
  output ex_ar_chan_Pop_mioi_wen_comp;
  output [67:0] ex_ar_chan_Pop_mioi_idat_mxwt;


  // Interconnect Declarations
  wire ex_ar_chan_Pop_mioi_biwt;
  wire ex_ar_chan_Pop_mioi_bdwt;
  wire [75:0] ex_ar_chan_Pop_mioi_idat;
  wire ex_ar_chan_Pop_mioi_irdy_ex_ar_process_sct;
  wire ex_ar_chan_Pop_mioi_ivld;
  wire [67:0] ex_ar_chan_Pop_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_conn_in_wait_v1 #(.width(32'sd76),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ex_ar_chan_Pop_mioi (
      .vld(ex_ar_chan_vld),
      .rdy(ex_ar_chan_rdy),
      .dat(ex_ar_chan_dat),
      .idat(ex_ar_chan_Pop_mioi_idat),
      .irdy(ex_ar_chan_Pop_mioi_irdy_ex_ar_process_sct),
      .ivld(ex_ar_chan_Pop_mioi_ivld),
      .clk(clk),
      .en(1'b0),
      .arst(rst_bar),
      .srst(1'b1)
    );
  axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_ex_ar_chan_Pop_mio_wait_ctrl
      axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_ex_ar_chan_Pop_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_ar_process_wen(ex_ar_process_wen),
      .ex_ar_process_wten(ex_ar_process_wten),
      .ex_ar_chan_Pop_mioi_oswt_unreg(ex_ar_chan_Pop_mioi_oswt_unreg),
      .ex_ar_chan_Pop_mioi_iswt0(ex_ar_chan_Pop_mioi_iswt0),
      .ex_ar_chan_Pop_mioi_biwt(ex_ar_chan_Pop_mioi_biwt),
      .ex_ar_chan_Pop_mioi_bdwt(ex_ar_chan_Pop_mioi_bdwt),
      .ex_ar_chan_Pop_mioi_irdy_ex_ar_process_sct(ex_ar_chan_Pop_mioi_irdy_ex_ar_process_sct),
      .ex_ar_chan_Pop_mioi_ivld(ex_ar_chan_Pop_mioi_ivld)
    );
  axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_ex_ar_chan_Pop_mio_wait_dp
      axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_ex_ar_chan_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_ar_chan_Pop_mioi_oswt_unreg(ex_ar_chan_Pop_mioi_oswt_unreg),
      .ex_ar_chan_Pop_mioi_bawt(ex_ar_chan_Pop_mioi_bawt),
      .ex_ar_chan_Pop_mioi_wen_comp(ex_ar_chan_Pop_mioi_wen_comp),
      .ex_ar_chan_Pop_mioi_idat_mxwt(ex_ar_chan_Pop_mioi_idat_mxwt_pconst),
      .ex_ar_chan_Pop_mioi_biwt(ex_ar_chan_Pop_mioi_biwt),
      .ex_ar_chan_Pop_mioi_bdwt(ex_ar_chan_Pop_mioi_bdwt),
      .ex_ar_chan_Pop_mioi_idat(ex_ar_chan_Pop_mioi_idat)
    );
  assign ex_ar_chan_Pop_mioi_idat_mxwt = ex_ar_chan_Pop_mioi_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_master_process
// ------------------------------------------------------------------


module scatter_gather_dma_master_process (
  clk, rst_bar, r_master0_r_vld, r_master0_r_rdy, r_master0_r_dat, dma_done_vld,
      dma_done_rdy, dma_done_dat, dma_cmd_chan_vld, dma_cmd_chan_rdy, dma_cmd_chan_dat,
      w_segment0_ex_aw_chan_vld, w_segment0_ex_aw_chan_rdy, w_segment0_ex_aw_chan_dat,
      w_segment0_w_chan_vld, w_segment0_w_chan_rdy, w_segment0_w_chan_dat, w_segment0_b_chan_vld,
      w_segment0_b_chan_rdy, w_segment0_b_chan_dat, r_segment0_ex_ar_chan_vld, r_segment0_ex_ar_chan_rdy,
      r_segment0_ex_ar_chan_dat
);
  input clk;
  input rst_bar;
  input r_master0_r_vld;
  output r_master0_r_rdy;
  input [70:0] r_master0_r_dat;
  output dma_done_vld;
  input dma_done_rdy;
  output dma_done_dat;
  input dma_cmd_chan_vld;
  output dma_cmd_chan_rdy;
  input [175:0] dma_cmd_chan_dat;
  output w_segment0_ex_aw_chan_vld;
  input w_segment0_ex_aw_chan_rdy;
  output [75:0] w_segment0_ex_aw_chan_dat;
  output w_segment0_w_chan_vld;
  input w_segment0_w_chan_rdy;
  output [72:0] w_segment0_w_chan_dat;
  input w_segment0_b_chan_vld;
  output w_segment0_b_chan_rdy;
  input [5:0] w_segment0_b_chan_dat;
  output r_segment0_ex_ar_chan_vld;
  input r_segment0_ex_ar_chan_rdy;
  output [75:0] r_segment0_ex_ar_chan_dat;


  // Interconnect Declarations
  wire master_process_wen;
  wire master_process_wten;
  wire dma_cmd_chan_Pop_mioi_wen_comp;
  wire [31:0] dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt;
  wire [31:0] dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt;
  wire [31:0] dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt;
  wire [31:0] dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt;
  wire [15:0] dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt;
  wire [15:0] dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt;
  wire r_segment0_ex_ar_chan_Push_mioi_wen_comp;
  wire w_segment0_ex_aw_chan_Push_mioi_wen_comp;
  wire r_master0_r_Pop_mioi_bawt;
  reg r_master0_r_Pop_mioi_iswt0;
  wire r_master0_r_Pop_mioi_wen_comp;
  wire [63:0] r_master0_r_Pop_mioi_idat_mxwt;
  wire w_segment0_w_chan_Push_mioi_bawt;
  wire w_segment0_w_chan_Push_mioi_wen_comp;
  reg [63:0] w_segment0_w_chan_Push_mioi_m_data_rsc_dat;
  wire w_segment0_b_chan_Pop_mioi_wen_comp;
  wire [1:0] w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt;
  wire dma_done_Push_mioi_wen_comp;
  reg dma_done_Push_mioi_idat_master_process;
  wire [16:0] fsm_output;
  wire operator_32_false_1_operator_32_false_1_nor_tmp;
  wire operator_32_false_4_operator_32_false_4_nor_tmp;
  wire and_dcpl_1;
  wire and_dcpl_5;
  wire and_dcpl_13;
  wire and_dcpl_30;
  wire and_dcpl_34;
  wire and_dcpl_42;
  wire or_dcpl_16;
  wire and_dcpl_47;
  wire or_dcpl_32;
  wire and_dcpl_60;
  wire or_dcpl_41;
  wire or_dcpl_45;
  wire or_dcpl_53;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_96;
  wire and_dcpl_99;
  wire and_dcpl_102;
  wire and_dcpl_105;
  wire or_dcpl_58;
  wire or_dcpl_61;
  wire or_dcpl_63;
  wire and_dcpl_107;
  wire and_dcpl_109;
  wire and_dcpl_112;
  wire and_dcpl_115;
  wire and_dcpl_118;
  wire or_dcpl_75;
  wire or_dcpl_80;
  wire and_dcpl_141;
  wire not_tmp_110;
  wire and_dcpl_145;
  wire and_tmp_7;
  wire and_dcpl_161;
  wire or_dcpl_96;
  wire and_dcpl_169;
  wire and_dcpl_184;
  wire or_tmp_122;
  wire or_tmp_135;
  wire or_tmp_147;
  wire or_tmp_173;
  wire and_336_cse;
  wire and_345_cse;
  wire and_390_cse;
  wire and_334_cse;
  wire and_335_cse;
  wire and_307_cse;
  reg while_case_0_while_stage_v;
  reg while_case_0_while_stage_0_1;
  reg while_case_1_while_while_stage_0_1;
  reg while_case_0_while_stage_v_1;
  reg while_case_2_while_while_stage_0_1;
  reg [15:0] while_cmd_dma_mode_sw_15_0_sva_st;
  reg while_case_1_while_while_stage_0;
  reg while_case_2_while_while_stage_0;
  reg while_case_0_while_stage_0;
  wire or_278_ssc;
  wire ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_mux_cse;
  wire ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_mux_1_cse;
  wire ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_1_mux_cse;
  wire ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_1_mux_1_cse;
  wire ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_2_mux_cse;
  wire ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_2_mux_1_cse;
  reg reg_dma_done_Push_mioi_iswt0_cse;
  reg reg_w_segment0_b_chan_Pop_mioi_iswt0_cse;
  reg reg_w_segment0_ex_aw_chan_Push_mioi_iswt0_cse;
  reg reg_r_segment0_ex_ar_chan_Push_mioi_iswt0_cse;
  reg reg_dma_cmd_chan_Pop_mioi_iswt0_cse;
  reg reg_w_segment0_w_chan_Push_mioi_iswt0_cse;
  wire or_89_cse;
  wire or_91_cse;
  wire or_93_cse;
  wire or_348_cse;
  wire and_639_cse;
  wire and_114_cse;
  wire or_198_rmff;
  reg master_process_flen_reg;
  wire and_rmff;
  wire or_203_rmff;
  wire or_201_rmff;
  wire [63:0] while_case_0_while_mux1h_2_rmff;
  wire or_193_rmff;
  reg [13:0] while_case_1_aw_ex_len_sva_13_0;
  wire or_tmp;
  wire [31:0] z_out;
  reg [31:0] while_cmd_total_len_sva;
  reg [31:0] while_cmd_scatter_stride_sva;
  reg [15:0] while_cmd_scatter_len_sva;
  reg [13:0] operator_17_true_2_acc_cse_sva;
  wire [14:0] nl_operator_17_true_2_acc_cse_sva;
  reg operator_32_false_1_slc_while_case_1_while_while_asn_incr_31_itm;
  reg operator_32_false_1_slc_while_case_1_while_while_asn_incr_29_itm;
  reg operator_32_false_1_slc_while_case_1_while_while_asn_incr_27_itm;
  reg operator_32_false_1_slc_while_case_1_while_while_asn_incr_23_itm;
  reg operator_32_false_1_slc_while_case_1_while_while_asn_incr_22_itm;
  reg operator_32_false_1_slc_while_case_1_while_while_asn_incr_15_itm;
  reg operator_32_false_1_slc_while_case_1_while_while_asn_incr_14_itm;
  reg operator_32_false_1_slc_while_case_1_while_while_asn_incr_13_itm;
  reg [31:0] while_case_1_while_acc_itm;
  wire while_case_0_while_stage_en_1_mx0w1;
  wire while_case_1_while_while_stage_en_2_mx0w1;
  wire while_case_1_while_while_stage_en_1_mx0w1;
  wire while_case_2_while_while_stage_en_1_mx0w1;
  wire [18:0] while_case_1_aw_ex_len_lpi_3_mx0_31_13;
  wire [18:0] while_case_2_ar_ex_len_lpi_3_mx0_31_13;
  wire [14:0] while_case_0_ar_ex_len_sva_mx3_27_13;
  wire or_168_tmp;
  wire or_267_rgt;
  wire while_case_0_ar_ex_len_and_rgt;
  wire and_255_rgt;
  wire while_case_0_ar_ex_len_and_2_rgt;
  wire or_276_rgt;
  wire operator_32_false_1_or_28_rgt;
  wire operator_32_false_1_or_30_rgt;
  wire operator_32_false_1_or_31_rgt;
  wire operator_32_false_1_and_49_rgt;
  wire while_case_0_ar_ex_len_and_4_ssc;
  reg [1:0] reg_while_case_0_ar_ex_len_ftd;
  reg [29:0] reg_while_case_0_ar_ex_len_ftd_1;
  wire while_cmd_scatter_len_and_cse;
  wire operator_32_false_1_and_53_cse;

  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_prb;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_1;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_1;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_2;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_2;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_3;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_3;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_4;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_4;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_5;
  wire ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_5;
  wire while_case_0_while_or_1_nl;
  wire mux1h_nl;
  wire nor_nl;
  wire while_case_0_while_mux_2_nl;
  wire while_case_0_while_mux_3_nl;
  wire nor_1_nl;
  wire while_case_1_while_while_mux_nl;
  wire while_case_1_while_while_mux_1_nl;
  wire nor_2_nl;
  wire while_case_2_while_while_mux_nl;
  wire while_case_2_while_while_mux_1_nl;
  wire or_205_nl;
  wire or_207_nl;
  wire or_208_nl;
  wire or_209_nl;
  wire while_switch_lp_mux_nl;
  wire or_232_nl;
  wire mux_29_nl;
  wire and_231_nl;
  wire while_switch_lp_mux1h_9_nl;
  wire and_405_nl;
  wire or_240_nl;
  wire mux_30_nl;
  wire while_case_1_while_while_mux_2_nl;
  wire while_case_1_while_while_mux1h_3_nl;
  wire nand_18_nl;
  wire mux_32_nl;
  wire nor_21_nl;
  wire and_435_nl;
  wire while_case_2_while_while_mux_2_nl;
  wire while_case_2_while_while_mux1h_3_nl;
  wire nand_17_nl;
  wire mux_34_nl;
  wire nor_20_nl;
  wire and_462_nl;
  wire while_case_0_ar_ex_len_and_5_nl;
  wire or_356_nl;
  wire while_case_0_while_mux1h_9_nl;
  wire while_switch_lp_while_switch_lp_or_4_nl;
  wire while_switch_lp_while_switch_lp_or_5_nl;
  wire while_switch_lp_while_switch_lp_or_6_nl;
  wire while_case_0_while_mux1h_14_nl;
  wire while_case_0_while_nor_1_nl;
  wire while_case_0_while_nor_2_nl;
  wire while_case_0_while_nor_3_nl;
  wire operator_32_false_1_and_48_nl;
  wire operator_32_false_1_and_52_nl;
  wire and_620_nl;
  wire and_622_nl;
  wire and_628_nl;
  wire and_630_nl;
  wire[32:0] acc_nl;
  wire[33:0] nl_acc_nl;
  wire[31:0] while_case_1_while_mux1h_2_nl;
  wire while_case_1_while_or_3_nl;
  wire while_case_1_while_or_4_nl;
  wire[31:0] while_case_1_while_while_case_1_while_or_1_nl;
  wire[31:0] while_case_1_while_mux_1_nl;
  wire while_case_1_while_or_5_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_inst_dma_cmd_chan_Pop_mioi_oswt_pff;
  assign nl_scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_inst_dma_cmd_chan_Pop_mioi_oswt_pff
      = fsm_output[1];
  wire [31:0] nl_scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_inst_r_segment0_ex_ar_chan_Push_mioi_m_addr_rsc_dat_master_process;
  assign nl_scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_inst_r_segment0_ex_ar_chan_Push_mioi_m_addr_rsc_dat_master_process
      = MUX_v_32_2_2(dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt, ({reg_while_case_0_ar_ex_len_ftd
      , reg_while_case_0_ar_ex_len_ftd_1}), fsm_output[10]);
  wire[29:0] while_switch_lp_while_switch_lp_mux_nl;
  wire [31:0] nl_scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_inst_r_segment0_ex_ar_chan_Push_mioi_m_ex_len_rsc_dat_master_process;
  assign while_switch_lp_while_switch_lp_mux_nl = MUX_v_30_2_2((z_out[29:0]), ({{16{while_case_1_aw_ex_len_sva_13_0[13]}},
      while_case_1_aw_ex_len_sva_13_0}), fsm_output[10]);
  assign nl_scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_inst_r_segment0_ex_ar_chan_Push_mioi_m_ex_len_rsc_dat_master_process
      = signext_32_30(while_switch_lp_while_switch_lp_mux_nl);
  wire [31:0] nl_scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_inst_w_segment0_ex_aw_chan_Push_mioi_m_addr_rsc_dat_master_process;
  assign nl_scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_inst_w_segment0_ex_aw_chan_Push_mioi_m_addr_rsc_dat_master_process
      = MUX_v_32_2_2(dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt, ({reg_while_case_0_ar_ex_len_ftd
      , reg_while_case_0_ar_ex_len_ftd_1}), fsm_output[5]);
  wire[29:0] while_switch_lp_while_switch_lp_mux_1_nl;
  wire [31:0] nl_scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_inst_w_segment0_ex_aw_chan_Push_mioi_m_ex_len_rsc_dat_master_process;
  assign while_switch_lp_while_switch_lp_mux_1_nl = MUX_v_30_2_2((z_out[29:0]), ({{16{while_case_1_aw_ex_len_sva_13_0[13]}},
      while_case_1_aw_ex_len_sva_13_0}), fsm_output[5]);
  assign nl_scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_inst_w_segment0_ex_aw_chan_Push_mioi_m_ex_len_rsc_dat_master_process
      = signext_32_30(while_switch_lp_while_switch_lp_mux_1_nl);
  wire  nl_scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_inst_w_segment0_w_chan_Push_mioi_oswt_unreg;
  assign nl_scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_inst_w_segment0_w_chan_Push_mioi_oswt_unreg
      = and_dcpl_60 & or_dcpl_80;
  wire  nl_scatter_gather_dma_master_process_master_process_fsm_inst_while_C_2_tr0;
  assign nl_scatter_gather_dma_master_process_master_process_fsm_inst_while_C_2_tr0
      = or_dcpl_53 | or_dcpl_45 | or_dcpl_41 | ((while_cmd_dma_mode_sw_15_0_sva_st[1:0]==2'b11));
  wire  nl_scatter_gather_dma_master_process_master_process_fsm_inst_while_C_2_tr1;
  assign nl_scatter_gather_dma_master_process_master_process_fsm_inst_while_C_2_tr1
      = and_dcpl_47;
  wire  nl_scatter_gather_dma_master_process_master_process_fsm_inst_while_C_2_tr2;
  assign nl_scatter_gather_dma_master_process_master_process_fsm_inst_while_C_2_tr2
      = and_dcpl_42 & and_dcpl_34 & and_dcpl_30 & (while_cmd_dma_mode_sw_15_0_sva_st[1:0]==2'b01);
  scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .dma_cmd_chan_vld(dma_cmd_chan_vld),
      .dma_cmd_chan_rdy(dma_cmd_chan_rdy),
      .dma_cmd_chan_dat(dma_cmd_chan_dat),
      .master_process_wen(master_process_wen),
      .dma_cmd_chan_Pop_mioi_oswt(reg_dma_cmd_chan_Pop_mioi_iswt0_cse),
      .dma_cmd_chan_Pop_mioi_wen_comp(dma_cmd_chan_Pop_mioi_wen_comp),
      .dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt(dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt),
      .dma_cmd_chan_Pop_mioi_oswt_pff(nl_scatter_gather_dma_master_process_dma_cmd_chan_Pop_mioi_inst_dma_cmd_chan_Pop_mioi_oswt_pff)
    );
  scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .r_segment0_ex_ar_chan_vld(r_segment0_ex_ar_chan_vld),
      .r_segment0_ex_ar_chan_rdy(r_segment0_ex_ar_chan_rdy),
      .r_segment0_ex_ar_chan_dat(r_segment0_ex_ar_chan_dat),
      .master_process_wen(master_process_wen),
      .r_segment0_ex_ar_chan_Push_mioi_oswt(reg_r_segment0_ex_ar_chan_Push_mioi_iswt0_cse),
      .r_segment0_ex_ar_chan_Push_mioi_wen_comp(r_segment0_ex_ar_chan_Push_mioi_wen_comp),
      .r_segment0_ex_ar_chan_Push_mioi_m_addr_rsc_dat_master_process(nl_scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_inst_r_segment0_ex_ar_chan_Push_mioi_m_addr_rsc_dat_master_process[31:0]),
      .r_segment0_ex_ar_chan_Push_mioi_m_ex_len_rsc_dat_master_process(nl_scatter_gather_dma_master_process_r_segment0_ex_ar_chan_Push_mioi_inst_r_segment0_ex_ar_chan_Push_mioi_m_ex_len_rsc_dat_master_process[31:0]),
      .r_segment0_ex_ar_chan_Push_mioi_oswt_pff(or_203_rmff)
    );
  scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_segment0_ex_aw_chan_vld(w_segment0_ex_aw_chan_vld),
      .w_segment0_ex_aw_chan_rdy(w_segment0_ex_aw_chan_rdy),
      .w_segment0_ex_aw_chan_dat(w_segment0_ex_aw_chan_dat),
      .master_process_wen(master_process_wen),
      .w_segment0_ex_aw_chan_Push_mioi_oswt(reg_w_segment0_ex_aw_chan_Push_mioi_iswt0_cse),
      .w_segment0_ex_aw_chan_Push_mioi_wen_comp(w_segment0_ex_aw_chan_Push_mioi_wen_comp),
      .w_segment0_ex_aw_chan_Push_mioi_m_addr_rsc_dat_master_process(nl_scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_inst_w_segment0_ex_aw_chan_Push_mioi_m_addr_rsc_dat_master_process[31:0]),
      .w_segment0_ex_aw_chan_Push_mioi_m_ex_len_rsc_dat_master_process(nl_scatter_gather_dma_master_process_w_segment0_ex_aw_chan_Push_mioi_inst_w_segment0_ex_aw_chan_Push_mioi_m_ex_len_rsc_dat_master_process[31:0]),
      .w_segment0_ex_aw_chan_Push_mioi_oswt_pff(or_201_rmff)
    );
  scatter_gather_dma_master_process_r_master0_r_Pop_mioi scatter_gather_dma_master_process_r_master0_r_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .r_master0_r_vld(r_master0_r_vld),
      .r_master0_r_rdy(r_master0_r_rdy),
      .r_master0_r_dat(r_master0_r_dat),
      .r_master0_r_Pop_mioi_oswt_unreg(or_198_rmff),
      .master_process_wen(master_process_wen),
      .master_process_wten(master_process_wten),
      .r_master0_r_Pop_mioi_bawt(r_master0_r_Pop_mioi_bawt),
      .r_master0_r_Pop_mioi_iswt0(r_master0_r_Pop_mioi_iswt0),
      .r_master0_r_Pop_mioi_wen_comp(r_master0_r_Pop_mioi_wen_comp),
      .r_master0_r_Pop_mioi_idat_mxwt(r_master0_r_Pop_mioi_idat_mxwt)
    );
  scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_segment0_w_chan_vld(w_segment0_w_chan_vld),
      .w_segment0_w_chan_rdy(w_segment0_w_chan_rdy),
      .w_segment0_w_chan_dat(w_segment0_w_chan_dat),
      .w_segment0_w_chan_Push_mioi_oswt_unreg(nl_scatter_gather_dma_master_process_w_segment0_w_chan_Push_mioi_inst_w_segment0_w_chan_Push_mioi_oswt_unreg),
      .master_process_wen(master_process_wen),
      .master_process_wten(master_process_wten),
      .w_segment0_w_chan_Push_mioi_bawt(w_segment0_w_chan_Push_mioi_bawt),
      .w_segment0_w_chan_Push_mioi_iswt0(reg_w_segment0_w_chan_Push_mioi_iswt0_cse),
      .w_segment0_w_chan_Push_mioi_wen_comp(w_segment0_w_chan_Push_mioi_wen_comp),
      .w_segment0_w_chan_Push_mioi_m_data_rsc_dat(while_case_0_while_mux1h_2_rmff),
      .w_segment0_w_chan_Push_mioi_iswt0_pff(or_198_rmff)
    );
  scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi scatter_gather_dma_master_process_w_segment0_b_chan_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_segment0_b_chan_vld(w_segment0_b_chan_vld),
      .w_segment0_b_chan_rdy(w_segment0_b_chan_rdy),
      .w_segment0_b_chan_dat(w_segment0_b_chan_dat),
      .master_process_wen(master_process_wen),
      .w_segment0_b_chan_Pop_mioi_oswt(reg_w_segment0_b_chan_Pop_mioi_iswt0_cse),
      .w_segment0_b_chan_Pop_mioi_wen_comp(w_segment0_b_chan_Pop_mioi_wen_comp),
      .w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt(w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt),
      .w_segment0_b_chan_Pop_mioi_oswt_pff(or_193_rmff)
    );
  scatter_gather_dma_master_process_dma_done_Push_mioi scatter_gather_dma_master_process_dma_done_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .dma_done_vld(dma_done_vld),
      .dma_done_rdy(dma_done_rdy),
      .dma_done_dat(dma_done_dat),
      .master_process_wen(master_process_wen),
      .dma_done_Push_mioi_oswt(reg_dma_done_Push_mioi_iswt0_cse),
      .dma_done_Push_mioi_wen_comp(dma_done_Push_mioi_wen_comp),
      .dma_done_Push_mioi_idat_master_process(dma_done_Push_mioi_idat_master_process)
    );
  scatter_gather_dma_master_process_staller_1 scatter_gather_dma_master_process_staller_1_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .master_process_flen_unreg(and_rmff),
      .master_process_wen(master_process_wen),
      .master_process_wten(master_process_wten),
      .dma_cmd_chan_Pop_mioi_wen_comp(dma_cmd_chan_Pop_mioi_wen_comp),
      .r_segment0_ex_ar_chan_Push_mioi_wen_comp(r_segment0_ex_ar_chan_Push_mioi_wen_comp),
      .w_segment0_ex_aw_chan_Push_mioi_wen_comp(w_segment0_ex_aw_chan_Push_mioi_wen_comp),
      .r_master0_r_Pop_mioi_wen_comp(r_master0_r_Pop_mioi_wen_comp),
      .w_segment0_w_chan_Push_mioi_wen_comp(w_segment0_w_chan_Push_mioi_wen_comp),
      .w_segment0_b_chan_Pop_mioi_wen_comp(w_segment0_b_chan_Pop_mioi_wen_comp),
      .dma_done_Push_mioi_wen_comp(dma_done_Push_mioi_wen_comp)
    );
  scatter_gather_dma_master_process_master_process_fsm scatter_gather_dma_master_process_master_process_fsm_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .master_process_wen(master_process_wen),
      .fsm_output(fsm_output),
      .while_C_2_tr0(nl_scatter_gather_dma_master_process_master_process_fsm_inst_while_C_2_tr0),
      .while_C_2_tr1(nl_scatter_gather_dma_master_process_master_process_fsm_inst_while_C_2_tr1),
      .while_C_2_tr2(nl_scatter_gather_dma_master_process_master_process_fsm_inst_while_C_2_tr2),
      .while_case_0_while_C_0_tr0(and_dcpl_92),
      .while_case_1_while_while_C_0_tr0(and_dcpl_94),
      .while_case_1_while_C_3_tr0(while_case_0_while_stage_v),
      .while_case_2_while_while_C_0_tr0(and_dcpl_96),
      .while_case_2_while_C_2_tr0(operator_32_false_4_operator_32_false_4_nor_tmp)
    );
  assign ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_mux_cse = MUX1HOT_s_1_1_2(1'b1,
      or_89_cse);
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_prb = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_mux_cse;
  // assert(true && "EmptyField should never be assigned or accessed") - /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/shared/pkgs/matchlib/cmod/include/UIntOrEmpty.h: line 38
  // psl default clock = (posedge clk);
  // psl scatter_gather_dma_master_process_UIntOrEmpty_h_ln38_assert_true_and_EmptyFieldshouldneverbeassignedoraccessed : assert always (  ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb  -> ptrue_EmptyField_should_never_be_assigned_or_accessed_prb );
  assign ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_mux_1_cse = MUX1HOT_s_1_1_2(master_process_wen,
      or_89_cse);
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_mux_1_cse;
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_1 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_mux_cse;
  // assert(true && "EmptyField should never be assigned or accessed") - /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/shared/pkgs/matchlib/cmod/include/UIntOrEmpty.h: line 38
  // psl scatter_gather_dma_master_process_UIntOrEmpty_h_ln38_assert_true_and_EmptyFieldshouldneverbeassignedoraccessed_1 : assert always (  ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_1  -> ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_1 );
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_1 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_mux_1_cse;
  assign ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_1_mux_cse = MUX1HOT_s_1_1_2(1'b1,
      or_91_cse);
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_2 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_1_mux_cse;
  // assert(true && "EmptyField should never be assigned or accessed") - /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/shared/pkgs/matchlib/cmod/include/UIntOrEmpty.h: line 38
  // psl scatter_gather_dma_master_process_UIntOrEmpty_h_ln38_assert_true_and_EmptyFieldshouldneverbeassignedoraccessed_2 : assert always (  ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_2  -> ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_2 );
  assign ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_1_mux_1_cse = MUX1HOT_s_1_1_2(master_process_wen,
      or_91_cse);
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_2 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_1_mux_1_cse;
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_3 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_1_mux_cse;
  // assert(true && "EmptyField should never be assigned or accessed") - /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/shared/pkgs/matchlib/cmod/include/UIntOrEmpty.h: line 38
  // psl scatter_gather_dma_master_process_UIntOrEmpty_h_ln38_assert_true_and_EmptyFieldshouldneverbeassignedoraccessed_3 : assert always (  ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_3  -> ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_3 );
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_3 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_1_mux_1_cse;
  assign ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_2_mux_cse = MUX1HOT_s_1_1_2(1'b1,
      or_93_cse);
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_4 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_2_mux_cse;
  // assert(true && "EmptyField should never be assigned or accessed") - /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/shared/pkgs/matchlib/cmod/include/UIntOrEmpty.h: line 38
  // psl scatter_gather_dma_master_process_UIntOrEmpty_h_ln38_assert_true_and_EmptyFieldshouldneverbeassignedoraccessed_4 : assert always (  ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_4  -> ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_4 );
  assign ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_2_mux_1_cse = MUX1HOT_s_1_1_2(master_process_wen,
      or_93_cse);
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_4 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_2_mux_1_cse;
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_5 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_2_mux_cse;
  // assert(true && "EmptyField should never be assigned or accessed") - /wv/hlsb/CATAPULT/10.6/PRODUCTION/aol/Mgc_home/shared/pkgs/matchlib/cmod/include/UIntOrEmpty.h: line 38
  // psl scatter_gather_dma_master_process_UIntOrEmpty_h_ln38_assert_true_and_EmptyFieldshouldneverbeassignedoraccessed_5 : assert always (  ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_5  -> ptrue_EmptyField_should_never_be_assigned_or_accessed_prb_5 );
  assign ptrue_EmptyField_should_never_be_assigned_or_accessed_ctrl_prb_5 = ar_burst_operator_enum_axi_AXI4_Encoding_AXBURST_unnamed_2_mux_1_cse;
  assign or_193_rmff = (and_dcpl_99 & (fsm_output[14])) | (fsm_output[8]);
  assign while_case_0_while_or_1_nl = (or_dcpl_61 & (fsm_output[7])) | (or_dcpl_63
      & (fsm_output[12])) | (~((fsm_output[12]) | (fsm_output[4]) | (fsm_output[7])))
      | and_307_cse;
  assign while_case_0_while_mux1h_2_rmff = MUX_v_64_2_2(r_master0_r_Pop_mioi_idat_mxwt,
      w_segment0_w_chan_Push_mioi_m_data_rsc_dat, while_case_0_while_or_1_nl);
  assign or_198_rmff = (and_dcpl_107 & (fsm_output[7])) | (and_dcpl_109 & (fsm_output[12]))
      | (and_dcpl_102 & (fsm_output[4]));
  assign or_201_rmff = (fsm_output[5]) | (and_dcpl_13 & and_dcpl_5 & and_dcpl_1 &
      (~ (dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[0])) & (fsm_output[2]));
  assign or_203_rmff = (fsm_output[10]) | (and_dcpl_13 & and_dcpl_5 & and_dcpl_1
      & (~ (dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[1])) & (fsm_output[2]));
  assign while_case_0_while_mux_2_nl = MUX_s_1_2_2(while_case_0_while_stage_0, while_case_0_while_stage_en_1_mx0w1,
      fsm_output[4]);
  assign while_case_0_while_mux_3_nl = MUX_s_1_2_2(while_case_0_while_stage_0_1,
      while_case_1_while_while_stage_en_2_mx0w1, fsm_output[4]);
  assign nor_nl = ~(((~(while_case_0_while_stage_v & (and_390_cse | and_307_cse)))
      & ((while_case_0_while_stage_0 & (~ or_tmp_122)) | (fsm_output[3]))) | while_case_0_while_mux_2_nl
      | while_case_0_while_mux_3_nl);
  assign while_case_1_while_while_mux_nl = MUX_s_1_2_2(while_case_1_while_while_stage_0,
      while_case_1_while_while_stage_en_1_mx0w1, fsm_output[7]);
  assign while_case_1_while_while_mux_1_nl = MUX_s_1_2_2(while_case_1_while_while_stage_0_1,
      while_case_1_while_while_stage_en_2_mx0w1, fsm_output[7]);
  assign nor_1_nl = ~(((~(while_case_0_while_stage_v & or_dcpl_61 & (fsm_output[7])))
      & ((while_case_1_while_while_stage_0 & (~ or_tmp_135)) | (fsm_output[6])))
      | while_case_1_while_while_mux_nl | while_case_1_while_while_mux_1_nl);
  assign while_case_2_while_while_mux_nl = MUX_s_1_2_2(while_case_2_while_while_stage_0,
      while_case_2_while_while_stage_en_1_mx0w1, fsm_output[12]);
  assign while_case_2_while_while_mux_1_nl = MUX_s_1_2_2(while_case_2_while_while_stage_0_1,
      while_case_1_while_while_stage_en_2_mx0w1, fsm_output[12]);
  assign nor_2_nl = ~(((~(while_case_0_while_stage_v & or_dcpl_63 & (fsm_output[12])))
      & ((while_case_2_while_while_stage_0 & (~ or_tmp_147)) | (fsm_output[11])))
      | while_case_2_while_while_mux_nl | while_case_2_while_while_mux_1_nl);
  assign or_205_nl = and_114_cse | ((or_dcpl_32 | while_case_0_while_stage_0 | while_case_0_while_stage_0_1)
      & (fsm_output[4]));
  assign or_207_nl = ((or_dcpl_32 | while_case_1_while_while_stage_0 | while_case_1_while_while_stage_0_1)
      & (fsm_output[7])) | (fsm_output[6]);
  assign or_208_nl = (fsm_output[11]) | ((or_dcpl_32 | while_case_2_while_while_stage_0
      | while_case_2_while_while_stage_0_1) & (fsm_output[12]));
  assign or_209_nl = (~((fsm_output[11]) | (fsm_output[6]) | (fsm_output[12]) | (fsm_output[4])
      | (fsm_output[7]) | (fsm_output[3]))) | and_345_cse;
  assign mux1h_nl = MUX1HOT_s_1_4_2(nor_nl, nor_1_nl, nor_2_nl, master_process_flen_reg,
      {or_205_nl , or_207_nl , or_208_nl , or_209_nl});
  assign and_rmff = mux1h_nl & (~(and_334_cse | and_335_cse | and_336_cse));
  assign or_267_rgt = (fsm_output[13]) | (fsm_output[8]);
  assign while_cmd_scatter_len_and_cse = master_process_wen & ((~ and_dcpl_161) |
      (fsm_output[0]) | (fsm_output[15]) | (fsm_output[14]) | (fsm_output[2]) | (fsm_output[4]));
  assign or_348_cse = (~ while_case_0_while_stage_v_1) | w_segment0_w_chan_Push_mioi_bawt;
  assign and_639_cse = or_348_cse & r_master0_r_Pop_mioi_bawt;
  assign or_168_tmp = and_dcpl_105 | or_dcpl_96;
  assign while_case_0_ar_ex_len_and_rgt = (dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[1])
      & (fsm_output[2]);
  assign and_255_rgt = (dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[1:0]==2'b01)
      & (fsm_output[2]);
  assign while_case_0_ar_ex_len_and_2_rgt = (~ or_168_tmp) & or_dcpl_80;
  assign or_276_rgt = (fsm_output[13]) | (fsm_output[9]);
  assign while_case_0_ar_ex_len_and_4_ssc = master_process_wen & (~(or_168_tmp &
      or_dcpl_80));
  assign and_114_cse = and_dcpl_47 & (fsm_output[3]);
  assign operator_32_false_1_or_28_rgt = (fsm_output[3]) | ((~ and_dcpl_184) & (fsm_output[4]));
  assign operator_32_false_1_or_30_rgt = (fsm_output[6]) | ((~ and_dcpl_184) & (fsm_output[7]));
  assign operator_32_false_1_or_31_rgt = (fsm_output[11]) | ((~ and_dcpl_184) & (fsm_output[12]));
  assign operator_32_false_1_and_53_cse = master_process_wen & (~((and_dcpl_184 &
      (fsm_output[4])) | (and_dcpl_184 & (fsm_output[7])) | (and_dcpl_184 & (fsm_output[12]))));
  assign operator_32_false_1_and_49_rgt = or_278_ssc & operator_32_false_1_or_28_rgt;
  assign or_89_cse = and_dcpl_13 & and_dcpl_5 & and_dcpl_1 & (dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[1:0]==2'b00)
      & (fsm_output[2]);
  assign or_91_cse = and_dcpl_13 & and_dcpl_5 & and_dcpl_1 & (dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[1:0]==2'b01)
      & (fsm_output[2]);
  assign or_93_cse = and_dcpl_13 & and_dcpl_5 & and_dcpl_1 & (dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[1:0]==2'b10)
      & (fsm_output[2]);
  assign while_case_0_while_stage_en_1_mx0w1 = while_case_0_while_stage_v & while_case_0_while_stage_0_1
      & r_master0_r_Pop_mioi_bawt & or_348_cse;
  assign while_case_1_while_while_stage_en_2_mx0w1 = while_case_0_while_stage_v_1
      & or_348_cse;
  assign while_case_1_while_while_stage_en_1_mx0w1 = while_case_0_while_stage_v &
      while_case_1_while_while_stage_0_1 & r_master0_r_Pop_mioi_bawt & or_348_cse;
  assign while_case_2_while_while_stage_en_1_mx0w1 = while_case_0_while_stage_v &
      while_case_2_while_while_stage_0_1 & r_master0_r_Pop_mioi_bawt & or_348_cse;
  assign while_case_0_ar_ex_len_sva_mx3_27_13 = MUX_v_15_2_2((reg_while_case_0_ar_ex_len_ftd_1[27:13]),
      (z_out[27:13]), or_278_ssc);
  assign operator_32_false_4_operator_32_false_4_nor_tmp = ~((z_out!=32'b00000000000000000000000000000000));
  assign and_620_nl = while_case_0_while_stage_v & (fsm_output[7]);
  assign and_622_nl = (~ while_case_0_while_stage_v) & (fsm_output[7]);
  assign while_case_1_aw_ex_len_lpi_3_mx0_31_13 = MUX1HOT_v_19_3_2((signext_19_1(while_case_1_aw_ex_len_sva_13_0[13])),
      (z_out[31:13]), ({reg_while_case_0_ar_ex_len_ftd , (reg_while_case_0_ar_ex_len_ftd_1[29:13])}),
      {(fsm_output[6]) , and_620_nl , and_622_nl});
  assign and_628_nl = while_case_0_while_stage_v & (fsm_output[12]);
  assign and_630_nl = (~ while_case_0_while_stage_v) & (fsm_output[12]);
  assign while_case_2_ar_ex_len_lpi_3_mx0_31_13 = MUX1HOT_v_19_3_2((signext_19_1(while_case_1_aw_ex_len_sva_13_0[13])),
      (z_out[31:13]), ({reg_while_case_0_ar_ex_len_ftd , (reg_while_case_0_ar_ex_len_ftd_1[29:13])}),
      {(fsm_output[11]) , and_628_nl , and_630_nl});
  assign operator_32_false_1_operator_32_false_1_nor_tmp = ~(operator_32_false_1_slc_while_case_1_while_while_asn_incr_31_itm
      | (reg_while_case_0_ar_ex_len_ftd[0]) | operator_32_false_1_slc_while_case_1_while_while_asn_incr_29_itm
      | (reg_while_case_0_ar_ex_len_ftd_1[28]) | operator_32_false_1_slc_while_case_1_while_while_asn_incr_27_itm
      | (reg_while_case_0_ar_ex_len_ftd_1[26:24]!=3'b000) | operator_32_false_1_slc_while_case_1_while_while_asn_incr_23_itm
      | operator_32_false_1_slc_while_case_1_while_while_asn_incr_22_itm | (reg_while_case_0_ar_ex_len_ftd_1[21:16]!=6'b000000)
      | operator_32_false_1_slc_while_case_1_while_while_asn_incr_15_itm | operator_32_false_1_slc_while_case_1_while_while_asn_incr_14_itm
      | operator_32_false_1_slc_while_case_1_while_while_asn_incr_13_itm | (reg_while_case_0_ar_ex_len_ftd_1[12:0]!=13'b0000000000000));
  assign and_dcpl_1 = ~((dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[15:14]!=2'b00));
  assign and_dcpl_5 = (dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[13:10]==4'b0000);
  assign and_dcpl_13 = (dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[9:2]==8'b00000000);
  assign and_dcpl_30 = ~((while_cmd_dma_mode_sw_15_0_sva_st[3:2]!=2'b00));
  assign and_dcpl_34 = (while_cmd_dma_mode_sw_15_0_sva_st[7:4]==4'b0000);
  assign and_dcpl_42 = (while_cmd_dma_mode_sw_15_0_sva_st[15:8]==8'b00000000);
  assign or_dcpl_16 = (fsm_output[11]) | (fsm_output[6]);
  assign and_dcpl_47 = and_dcpl_42 & and_dcpl_34 & and_dcpl_30 & (while_cmd_dma_mode_sw_15_0_sva_st[1:0]==2'b00);
  assign or_dcpl_32 = ~(while_case_0_while_stage_v_1 & w_segment0_w_chan_Push_mioi_bawt);
  assign and_dcpl_60 = while_case_0_while_stage_v_1 & w_segment0_w_chan_Push_mioi_bawt;
  assign or_dcpl_41 = (while_cmd_dma_mode_sw_15_0_sva_st[3:2]!=2'b00);
  assign or_dcpl_45 = (while_cmd_dma_mode_sw_15_0_sva_st[7:4]!=4'b0000);
  assign or_dcpl_53 = (while_cmd_dma_mode_sw_15_0_sva_st[15:8]!=8'b00000000);
  assign and_dcpl_92 = and_dcpl_60 & (~ while_case_0_while_stage_0) & (~ while_case_0_while_stage_0_1);
  assign and_dcpl_94 = and_dcpl_60 & (~ while_case_1_while_while_stage_0) & (~ while_case_1_while_while_stage_0_1);
  assign and_dcpl_96 = and_dcpl_60 & (~ while_case_2_while_while_stage_0) & (~ while_case_2_while_while_stage_0_1);
  assign and_dcpl_99 = and_dcpl_42 & and_dcpl_34 & and_dcpl_30 & (~ (while_cmd_dma_mode_sw_15_0_sva_st[0]));
  assign and_dcpl_102 = and_639_cse & while_case_0_while_stage_v & while_case_0_while_stage_0_1;
  assign and_dcpl_105 = while_case_0_while_stage_v_1 & (~ w_segment0_w_chan_Push_mioi_bawt);
  assign or_dcpl_58 = and_dcpl_105 | (~ r_master0_r_Pop_mioi_bawt);
  assign or_dcpl_61 = or_dcpl_58 | (~ while_case_0_while_stage_v) | (~ while_case_1_while_while_stage_0_1);
  assign or_dcpl_63 = or_dcpl_58 | (~ while_case_0_while_stage_v) | (~ while_case_2_while_while_stage_0_1);
  assign and_dcpl_107 = and_639_cse & while_case_0_while_stage_v & while_case_1_while_while_stage_0_1;
  assign and_dcpl_109 = and_639_cse & while_case_0_while_stage_v & while_case_2_while_while_stage_0_1;
  assign and_dcpl_112 = (~((~(and_639_cse & (~ operator_32_false_1_operator_32_false_1_nor_tmp)
      & while_case_1_while_while_stage_0_1)) & while_case_0_while_stage_v)) & while_case_1_while_while_stage_0;
  assign and_dcpl_115 = (~((~(and_639_cse & (~ operator_32_false_1_operator_32_false_1_nor_tmp)
      & while_case_2_while_while_stage_0_1)) & while_case_0_while_stage_v)) & while_case_2_while_while_stage_0;
  assign and_dcpl_118 = (~((~(and_639_cse & (~ operator_32_false_1_operator_32_false_1_nor_tmp)
      & while_case_0_while_stage_0_1)) & while_case_0_while_stage_v)) & while_case_0_while_stage_0;
  assign or_dcpl_75 = (while_cmd_dma_mode_sw_15_0_sva_st[1:0]!=2'b00);
  assign or_dcpl_80 = (fsm_output[12]) | (fsm_output[4]) | (fsm_output[7]);
  assign and_dcpl_141 = while_case_0_while_stage_v & operator_32_false_1_operator_32_false_1_nor_tmp;
  assign not_tmp_110 = ~(while_case_0_while_stage_0 | or_dcpl_32);
  assign and_dcpl_145 = while_case_0_while_stage_v & (~ operator_32_false_1_operator_32_false_1_nor_tmp);
  assign and_tmp_7 = while_case_0_while_stage_v & r_master0_r_Pop_mioi_bawt & or_348_cse;
  assign and_dcpl_161 = ~((fsm_output[16]) | (fsm_output[1]));
  assign or_dcpl_96 = ~(r_master0_r_Pop_mioi_bawt & while_case_0_while_stage_v);
  assign and_dcpl_169 = r_master0_r_Pop_mioi_bawt & while_case_0_while_stage_v;
  assign and_dcpl_184 = or_dcpl_58 & while_case_0_while_stage_v;
  assign and_307_cse = (or_dcpl_58 | (~ while_case_0_while_stage_v) | (~ while_case_0_while_stage_0_1))
      & (fsm_output[4]);
  assign and_336_cse = and_dcpl_92 & (fsm_output[4]);
  assign and_334_cse = and_dcpl_94 & (fsm_output[7]);
  assign and_335_cse = and_dcpl_96 & (fsm_output[12]);
  assign and_345_cse = (or_dcpl_53 | or_dcpl_45 | or_dcpl_41 | or_dcpl_75) & (fsm_output[3]);
  assign or_tmp_122 = and_639_cse & and_dcpl_141 & while_case_0_while_stage_0_1 &
      (fsm_output[4]);
  assign and_390_cse = ~((fsm_output[4:3]!=2'b00));
  assign or_tmp_135 = and_639_cse & and_dcpl_141 & while_case_1_while_while_stage_0_1
      & (fsm_output[7]);
  assign or_tmp_147 = and_639_cse & and_dcpl_141 & while_case_2_while_while_stage_0_1
      & (fsm_output[12]);
  assign or_tmp_173 = or_dcpl_16 | (fsm_output[3]);
  assign or_278_ssc = while_case_0_while_stage_v & (fsm_output[4]);
  assign or_tmp = (fsm_output[10]) | (fsm_output[5]);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      dma_done_Push_mioi_idat_master_process <= 1'b0;
      reg_dma_done_Push_mioi_iswt0_cse <= 1'b0;
      reg_w_segment0_b_chan_Pop_mioi_iswt0_cse <= 1'b0;
      w_segment0_w_chan_Push_mioi_m_data_rsc_dat <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      reg_w_segment0_w_chan_Push_mioi_iswt0_cse <= 1'b0;
      r_master0_r_Pop_mioi_iswt0 <= 1'b0;
      reg_w_segment0_ex_aw_chan_Push_mioi_iswt0_cse <= 1'b0;
      reg_r_segment0_ex_ar_chan_Push_mioi_iswt0_cse <= 1'b0;
      reg_dma_cmd_chan_Pop_mioi_iswt0_cse <= 1'b0;
      master_process_flen_reg <= 1'b0;
      while_case_0_while_stage_0 <= 1'b0;
      while_case_0_while_stage_0_1 <= 1'b0;
      while_case_1_while_while_stage_0 <= 1'b0;
      while_case_1_while_while_stage_0_1 <= 1'b0;
      while_case_2_while_while_stage_0 <= 1'b0;
      while_case_2_while_while_stage_0_1 <= 1'b0;
      while_case_0_while_stage_v <= 1'b0;
      while_case_0_while_stage_v_1 <= 1'b0;
    end
    else if ( master_process_wen ) begin
      dma_done_Push_mioi_idat_master_process <= ~((w_segment0_b_chan_Pop_mioi_return_resp_rsc_z_mxwt!=2'b00));
      reg_dma_done_Push_mioi_iswt0_cse <= (and_dcpl_99 & (fsm_output[15])) | (while_case_0_while_stage_v
          & (fsm_output[9]));
      reg_w_segment0_b_chan_Pop_mioi_iswt0_cse <= or_193_rmff;
      w_segment0_w_chan_Push_mioi_m_data_rsc_dat <= while_case_0_while_mux1h_2_rmff;
      reg_w_segment0_w_chan_Push_mioi_iswt0_cse <= or_198_rmff;
      r_master0_r_Pop_mioi_iswt0 <= (and_dcpl_112 & (fsm_output[7])) | or_dcpl_16
          | and_114_cse | (and_dcpl_115 & (fsm_output[12])) | (and_dcpl_118 & (fsm_output[4]));
      reg_w_segment0_ex_aw_chan_Push_mioi_iswt0_cse <= or_201_rmff;
      reg_r_segment0_ex_ar_chan_Push_mioi_iswt0_cse <= or_203_rmff;
      reg_dma_cmd_chan_Pop_mioi_iswt0_cse <= fsm_output[1];
      master_process_flen_reg <= and_rmff;
      while_case_0_while_stage_0 <= (while_switch_lp_mux_nl & (~ or_tmp_122)) | and_114_cse;
      while_case_0_while_stage_0_1 <= (while_switch_lp_mux1h_9_nl & (~ or_tmp_122))
          | and_114_cse;
      while_case_1_while_while_stage_0 <= (while_case_1_while_while_mux_2_nl & (~
          or_tmp_135)) | (fsm_output[6]);
      while_case_1_while_while_stage_0_1 <= (while_case_1_while_while_mux1h_3_nl
          & (~ or_tmp_135)) | (fsm_output[6]);
      while_case_2_while_while_stage_0 <= (while_case_2_while_while_mux_2_nl & (~
          or_tmp_147)) | (fsm_output[11]);
      while_case_2_while_while_stage_0_1 <= (while_case_2_while_while_mux1h_3_nl
          & (~ or_tmp_147)) | (fsm_output[11]);
      while_case_0_while_stage_v <= while_case_0_while_mux1h_9_nl | or_tmp_173;
      while_case_0_while_stage_v_1 <= ~(while_case_0_while_mux1h_14_nl | or_tmp_173);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_cmd_total_len_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( master_process_wen & (~((fsm_output[5]) | (fsm_output[10]) | or_dcpl_16
        | (fsm_output[9]) | (fsm_output[12]) | (fsm_output[7]) | (fsm_output[3])))
        ) begin
      while_cmd_total_len_sva <= MUX_v_32_2_2(dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt,
          z_out, or_267_rgt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_cmd_scatter_len_sva <= 16'b0000000000000000;
      operator_17_true_2_acc_cse_sva <= 14'b00000000000000;
      while_cmd_scatter_stride_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( while_cmd_scatter_len_and_cse ) begin
      while_cmd_scatter_len_sva <= dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt;
      operator_17_true_2_acc_cse_sva <= nl_operator_17_true_2_acc_cse_sva[13:0];
      while_cmd_scatter_stride_sva <= dma_cmd_chan_Pop_mioi_return_scatter_stride_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_cmd_dma_mode_sw_15_0_sva_st <= 16'b0000000000000000;
    end
    else if ( master_process_wen & ((~ and_dcpl_161) | (fsm_output[0]) | (fsm_output[15])
        | (fsm_output[2])) ) begin
      while_cmd_dma_mode_sw_15_0_sva_st <= dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      reg_while_case_0_ar_ex_len_ftd <= 2'b00;
    end
    else if ( while_case_0_ar_ex_len_and_4_ssc & (~(or_dcpl_75 & (fsm_output[3])))
        ) begin
      reg_while_case_0_ar_ex_len_ftd <= MUX1HOT_v_2_6_2((dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt[31:30]),
          (dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt[31:30]), (signext_2_1(reg_while_case_0_ar_ex_len_ftd_1[29])),
          (z_out[31:30]), (signext_2_1(while_case_1_aw_ex_len_sva_13_0[13])), (while_case_1_while_acc_itm[31:30]),
          {while_case_0_ar_ex_len_and_rgt , and_255_rgt , while_case_0_ar_ex_len_and_5_nl
          , while_case_0_ar_ex_len_and_2_rgt , or_dcpl_16 , or_276_rgt});
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      reg_while_case_0_ar_ex_len_ftd_1 <= 30'b000000000000000000000000000000;
    end
    else if ( while_case_0_ar_ex_len_and_4_ssc & (~ (fsm_output[3])) ) begin
      reg_while_case_0_ar_ex_len_ftd_1 <= MUX1HOT_v_30_5_2((dma_cmd_chan_Pop_mioi_return_ar_addr_rsc_z_mxwt[29:0]),
          (dma_cmd_chan_Pop_mioi_return_aw_addr_rsc_z_mxwt[29:0]), ({{16{while_case_1_aw_ex_len_sva_13_0[13]}},
          while_case_1_aw_ex_len_sva_13_0}), (while_case_1_while_acc_itm[29:0]),
          (z_out[29:0]), {while_case_0_ar_ex_len_and_rgt , and_255_rgt , or_dcpl_16
          , or_276_rgt , or_356_nl});
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_case_1_aw_ex_len_sva_13_0 <= 14'b00000000000000;
    end
    else if ( master_process_wen & ((fsm_output[13]) | (fsm_output[9]) | (fsm_output[3]))
        ) begin
      while_case_1_aw_ex_len_sva_13_0 <= operator_17_true_2_acc_cse_sva;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_13_itm <= 1'b0;
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_14_itm <= 1'b0;
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_15_itm <= 1'b0;
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_22_itm <= 1'b0;
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_23_itm <= 1'b0;
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_27_itm <= 1'b0;
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_29_itm <= 1'b0;
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_31_itm <= 1'b0;
    end
    else if ( operator_32_false_1_and_53_cse ) begin
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_13_itm <= MUX1HOT_s_1_3_2((while_case_0_ar_ex_len_sva_mx3_27_13[0]),
          (while_case_1_aw_ex_len_lpi_3_mx0_31_13[0]), (while_case_2_ar_ex_len_lpi_3_mx0_31_13[0]),
          {operator_32_false_1_or_28_rgt , operator_32_false_1_or_30_rgt , operator_32_false_1_or_31_rgt});
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_14_itm <= MUX1HOT_s_1_3_2((while_case_0_ar_ex_len_sva_mx3_27_13[1]),
          (while_case_1_aw_ex_len_lpi_3_mx0_31_13[1]), (while_case_2_ar_ex_len_lpi_3_mx0_31_13[1]),
          {operator_32_false_1_or_28_rgt , operator_32_false_1_or_30_rgt , operator_32_false_1_or_31_rgt});
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_15_itm <= MUX1HOT_s_1_3_2((while_case_0_ar_ex_len_sva_mx3_27_13[2]),
          (while_case_1_aw_ex_len_lpi_3_mx0_31_13[2]), (while_case_2_ar_ex_len_lpi_3_mx0_31_13[2]),
          {operator_32_false_1_or_28_rgt , operator_32_false_1_or_30_rgt , operator_32_false_1_or_31_rgt});
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_22_itm <= MUX1HOT_s_1_3_2((while_case_0_ar_ex_len_sva_mx3_27_13[9]),
          (while_case_1_aw_ex_len_lpi_3_mx0_31_13[9]), (while_case_2_ar_ex_len_lpi_3_mx0_31_13[9]),
          {operator_32_false_1_or_28_rgt , operator_32_false_1_or_30_rgt , operator_32_false_1_or_31_rgt});
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_23_itm <= MUX1HOT_s_1_3_2((while_case_0_ar_ex_len_sva_mx3_27_13[10]),
          (while_case_1_aw_ex_len_lpi_3_mx0_31_13[10]), (while_case_2_ar_ex_len_lpi_3_mx0_31_13[10]),
          {operator_32_false_1_or_28_rgt , operator_32_false_1_or_30_rgt , operator_32_false_1_or_31_rgt});
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_27_itm <= MUX1HOT_s_1_3_2((while_case_0_ar_ex_len_sva_mx3_27_13[14]),
          (while_case_1_aw_ex_len_lpi_3_mx0_31_13[14]), (while_case_2_ar_ex_len_lpi_3_mx0_31_13[14]),
          {operator_32_false_1_or_28_rgt , operator_32_false_1_or_30_rgt , operator_32_false_1_or_31_rgt});
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_29_itm <= MUX1HOT_s_1_4_2((reg_while_case_0_ar_ex_len_ftd_1[29]),
          (z_out[29]), (while_case_1_aw_ex_len_lpi_3_mx0_31_13[16]), (while_case_2_ar_ex_len_lpi_3_mx0_31_13[16]),
          {operator_32_false_1_and_48_nl , operator_32_false_1_and_49_rgt , operator_32_false_1_or_30_rgt
          , operator_32_false_1_or_31_rgt});
      operator_32_false_1_slc_while_case_1_while_while_asn_incr_31_itm <= MUX1HOT_s_1_5_2((reg_while_case_0_ar_ex_len_ftd_1[29]),
          (z_out[31]), (reg_while_case_0_ar_ex_len_ftd[1]), (while_case_1_aw_ex_len_lpi_3_mx0_31_13[18]),
          (while_case_2_ar_ex_len_lpi_3_mx0_31_13[18]), {(fsm_output[3]) , operator_32_false_1_and_49_rgt
          , operator_32_false_1_and_52_nl , operator_32_false_1_or_30_rgt , operator_32_false_1_or_31_rgt});
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_case_1_while_acc_itm <= 32'b00000000000000000000000000000000;
    end
    else if ( master_process_wen & (~(or_dcpl_16 | (fsm_output[8]) | (fsm_output[12])
        | (fsm_output[7]))) ) begin
      while_case_1_while_acc_itm <= z_out;
    end
  end
  assign and_231_nl = operator_32_false_1_operator_32_false_1_nor_tmp & while_case_0_while_stage_v
      & r_master0_r_Pop_mioi_bawt & or_348_cse;
  assign mux_29_nl = MUX_s_1_2_2(not_tmp_110, and_231_nl, while_case_0_while_stage_0_1);
  assign or_232_nl = and_390_cse | and_345_cse | ((~ mux_29_nl) & (fsm_output[4]));
  assign while_switch_lp_mux_nl = MUX_s_1_2_2(while_case_0_while_stage_en_1_mx0w1,
      while_case_0_while_stage_0, or_232_nl);
  assign and_405_nl = and_639_cse & and_dcpl_145 & while_case_0_while_stage_0_1 &
      (fsm_output[4]);
  assign mux_30_nl = MUX_s_1_2_2(not_tmp_110, and_tmp_7, while_case_0_while_stage_0_1);
  assign or_240_nl = and_390_cse | and_345_cse | ((~ mux_30_nl) & (fsm_output[4]));
  assign while_switch_lp_mux1h_9_nl = MUX1HOT_s_1_3_2(while_case_0_while_stage_0,
      while_case_1_while_while_stage_en_2_mx0w1, while_case_0_while_stage_0_1, {and_405_nl
      , and_336_cse , or_240_nl});
  assign while_case_1_while_while_mux_2_nl = MUX_s_1_2_2(while_case_1_while_while_stage_0,
      while_case_1_while_while_stage_en_1_mx0w1, and_334_cse);
  assign nor_21_nl = ~(while_case_1_while_while_stage_0 | or_dcpl_32);
  assign mux_32_nl = MUX_s_1_2_2(nor_21_nl, and_tmp_7, while_case_1_while_while_stage_0_1);
  assign nand_18_nl = ~((fsm_output[7]) & mux_32_nl);
  assign and_435_nl = and_639_cse & and_dcpl_145 & while_case_1_while_while_stage_0_1
      & (fsm_output[7]);
  assign while_case_1_while_while_mux1h_3_nl = MUX1HOT_s_1_3_2(while_case_1_while_while_stage_0_1,
      while_case_1_while_while_stage_0, while_case_1_while_while_stage_en_2_mx0w1,
      {nand_18_nl , and_435_nl , and_334_cse});
  assign while_case_2_while_while_mux_2_nl = MUX_s_1_2_2(while_case_2_while_while_stage_0,
      while_case_2_while_while_stage_en_1_mx0w1, and_335_cse);
  assign nor_20_nl = ~(while_case_2_while_while_stage_0 | or_dcpl_32);
  assign mux_34_nl = MUX_s_1_2_2(nor_20_nl, and_tmp_7, while_case_2_while_while_stage_0_1);
  assign nand_17_nl = ~((fsm_output[12]) & mux_34_nl);
  assign and_462_nl = and_639_cse & and_dcpl_145 & while_case_2_while_while_stage_0_1
      & (fsm_output[12]);
  assign while_case_2_while_while_mux1h_3_nl = MUX1HOT_s_1_3_2(while_case_2_while_while_stage_0_1,
      while_case_2_while_while_stage_0, while_case_1_while_while_stage_en_2_mx0w1,
      {nand_17_nl , and_462_nl , and_335_cse});
  assign while_switch_lp_while_switch_lp_or_4_nl = (while_case_0_while_stage_v &
      (~(or_348_cse & (operator_32_false_1_operator_32_false_1_nor_tmp | (~ while_case_0_while_stage_0))
      & and_dcpl_169 & while_case_0_while_stage_0_1))) | and_dcpl_118;
  assign while_switch_lp_while_switch_lp_or_5_nl = (while_case_0_while_stage_v &
      (~(or_348_cse & (operator_32_false_1_operator_32_false_1_nor_tmp | (~ while_case_1_while_while_stage_0))
      & and_dcpl_169 & while_case_1_while_while_stage_0_1))) | and_dcpl_112;
  assign while_switch_lp_while_switch_lp_or_6_nl = (while_case_0_while_stage_v &
      (~(or_348_cse & (operator_32_false_1_operator_32_false_1_nor_tmp | (~ while_case_2_while_while_stage_0))
      & and_dcpl_169 & while_case_2_while_while_stage_0_1))) | and_dcpl_115;
  assign while_case_0_while_mux1h_9_nl = MUX1HOT_s_1_4_2(while_switch_lp_while_switch_lp_or_4_nl,
      while_switch_lp_while_switch_lp_or_5_nl, operator_32_false_4_operator_32_false_4_nor_tmp,
      while_switch_lp_while_switch_lp_or_6_nl, {(fsm_output[4]) , (fsm_output[7])
      , (fsm_output[8]) , (fsm_output[12])});
  assign while_case_0_while_nor_1_nl = ~((while_case_0_while_stage_v_1 & (~((or_dcpl_96
      | (~ while_case_0_while_stage_0_1)) & and_dcpl_60))) | and_dcpl_102);
  assign while_case_0_while_nor_2_nl = ~((while_case_0_while_stage_v_1 & (~((or_dcpl_96
      | (~ while_case_1_while_while_stage_0_1)) & and_dcpl_60))) | and_dcpl_107);
  assign while_case_0_while_nor_3_nl = ~((while_case_0_while_stage_v_1 & (~((or_dcpl_96
      | (~ while_case_2_while_while_stage_0_1)) & and_dcpl_60))) | and_dcpl_109);
  assign while_case_0_while_mux1h_14_nl = MUX1HOT_s_1_3_2(while_case_0_while_nor_1_nl,
      while_case_0_while_nor_2_nl, while_case_0_while_nor_3_nl, {(fsm_output[4])
      , (fsm_output[7]) , (fsm_output[12])});
  assign nl_operator_17_true_2_acc_cse_sva  = conv_u2s_13_14(dma_cmd_chan_Pop_mioi_return_scatter_len_rsc_z_mxwt[15:3])
      + 14'b11111111111111;
  assign while_case_0_ar_ex_len_and_5_nl = (~ or_dcpl_75) & (fsm_output[3]);
  assign or_356_nl = ((dma_cmd_chan_Pop_mioi_return_dma_mode_rsc_z_mxwt[1:0]==2'b00)
      & (fsm_output[2])) | while_case_0_ar_ex_len_and_2_rgt;
  assign operator_32_false_1_and_48_nl = (~ or_278_ssc) & operator_32_false_1_or_28_rgt;
  assign operator_32_false_1_and_52_nl = (and_390_cse | ((~ while_case_0_while_stage_v)
      & (fsm_output[4]))) & operator_32_false_1_or_28_rgt;
  assign while_case_1_while_or_3_nl = or_tmp | or_dcpl_80;
  assign while_case_1_while_mux1h_2_nl = MUX1HOT_v_32_3_2(({reg_while_case_0_ar_ex_len_ftd
      , reg_while_case_0_ar_ex_len_ftd_1}), ({3'b000 , (dma_cmd_chan_Pop_mioi_return_total_len_rsc_z_mxwt[31:3])}),
      while_cmd_total_len_sva, {while_case_1_while_or_3_nl , (fsm_output[2]) , or_267_rgt});
  assign while_case_1_while_or_4_nl = (~(or_tmp | (fsm_output[2]) | or_dcpl_80))
      | or_267_rgt;
  assign while_case_1_while_mux_1_nl = MUX_v_32_2_2(while_cmd_scatter_stride_sva,
      ({16'b1111111111111111 , (~ while_cmd_scatter_len_sva)}), or_267_rgt);
  assign while_case_1_while_or_5_nl = (fsm_output[2]) | or_dcpl_80;
  assign while_case_1_while_while_case_1_while_or_1_nl = MUX_v_32_2_2(while_case_1_while_mux_1_nl,
      32'b11111111111111111111111111111111, while_case_1_while_or_5_nl);
  assign nl_acc_nl = ({while_case_1_while_mux1h_2_nl , while_case_1_while_or_4_nl})
      + ({while_case_1_while_while_case_1_while_or_1_nl , 1'b1});
  assign acc_nl = nl_acc_nl[32:0];
  assign z_out = readslicef_33_32_1(acc_nl);

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & {1{sel}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & {1{sel}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & {1{sel}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & {1{sel}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [18:0] MUX1HOT_v_19_3_2;
    input [18:0] input_2;
    input [18:0] input_1;
    input [18:0] input_0;
    input [2:0] sel;
    reg [18:0] result;
  begin
    result = input_0 & {19{sel[0]}};
    result = result | ( input_1 & {19{sel[1]}});
    result = result | ( input_2 & {19{sel[2]}});
    MUX1HOT_v_19_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_6_2;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [5:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    result = result | ( input_4 & {2{sel[4]}});
    result = result | ( input_5 & {2{sel[5]}});
    MUX1HOT_v_2_6_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_5_2;
    input [29:0] input_4;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [4:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    result = result | ( input_3 & {30{sel[3]}});
    result = result | ( input_4 & {30{sel[4]}});
    MUX1HOT_v_30_5_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input  sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input  sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [31:0] readslicef_33_32_1;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_33_32_1 = tmp[31:0];
  end
  endfunction


  function automatic [18:0] signext_19_1;
    input  vector;
  begin
    signext_19_1= {{18{vector}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [31:0] signext_32_30;
    input [29:0] vector;
  begin
    signext_32_30= {{2{vector[29]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_u2s_13_14 ;
    input [12:0]  vector ;
  begin
    conv_u2s_13_14 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma_slave_process
// ------------------------------------------------------------------


module scatter_gather_dma_slave_process (
  clk, rst_bar, w_slave0_aw_vld, w_slave0_aw_rdy, w_slave0_aw_dat, w_slave0_w_vld,
      w_slave0_w_rdy, w_slave0_w_dat, w_slave0_b_vld, w_slave0_b_rdy, w_slave0_b_dat,
      dma_cmd_chan_vld, dma_cmd_chan_rdy, dma_cmd_chan_dat
);
  input clk;
  input rst_bar;
  input w_slave0_aw_vld;
  output w_slave0_aw_rdy;
  input [31:0] w_slave0_aw_dat;
  input w_slave0_w_vld;
  output w_slave0_w_rdy;
  input [31:0] w_slave0_w_dat;
  output w_slave0_b_vld;
  input w_slave0_b_rdy;
  output [1:0] w_slave0_b_dat;
  output dma_cmd_chan_vld;
  input dma_cmd_chan_rdy;
  output [175:0] dma_cmd_chan_dat;


  // Interconnect Declarations
  wire slave_process_wen;
  wire w_slave0_aw_Pop_mioi_wen_comp;
  wire [31:0] w_slave0_aw_Pop_mioi_idat_mxwt;
  wire w_slave0_w_Pop_mioi_wen_comp;
  wire [31:0] w_slave0_w_Pop_mioi_idat_mxwt;
  wire dma_cmd_chan_Push_mioi_wen_comp;
  wire w_slave0_b_Push_mioi_wen_comp;
  reg w_slave0_b_Push_mioi_idat_slave_process_1;
  wire [2:0] fsm_output;
  wire while_case_28_if_1_oif_1_unequal_tmp;
  wire while_case_28_if_while_case_28_if_or_1_tmp;
  wire while_switch_lp_while_switch_lp_nor_1_tmp;
  wire while_switch_lp_nor_6_tmp;
  wire while_switch_lp_nor_5_tmp;
  wire while_switch_lp_nor_4_tmp;
  wire while_switch_lp_nor_3_tmp;
  wire while_switch_lp_nor_2_tmp;
  wire while_switch_lp_nor_1_tmp;
  wire or_dcpl_1;
  wire or_dcpl_5;
  wire or_dcpl_11;
  wire or_dcpl_17;
  wire or_dcpl_27;
  wire or_dcpl_31;
  wire and_dcpl_47;
  reg [31:0] cmd1_scatter_stride_sva;
  reg [15:0] cmd1_scatter_len_sva;
  wire while_switch_lp_equal_tmp_7;
  wire while_switch_lp_equal_tmp_8;
  wire while_switch_lp_equal_tmp_9;
  wire while_switch_lp_equal_tmp_10;
  wire while_switch_lp_equal_tmp_11;
  reg [15:0] cmd1_dma_mode_sva;
  reg while_case_28_if_1_lor_lpi_1_dfm;
  wire while_case_28_if_1_lor_lpi_1_dfm_mx0w0;
  reg reg_w_slave0_b_Push_mioi_iswt0_cse;
  reg reg_dma_cmd_chan_Push_mioi_iswt0_cse;
  reg reg_w_slave0_w_Pop_mioi_iswt0_cse;
  wire or_cse;
  wire and_72_cse;
  wire and_50_rmff;
  reg [31:0] cmd1_ar_addr_sva;
  reg [31:0] cmd1_aw_addr_sva;
  reg [31:0] cmd1_total_len_sva;
  reg [15:0] cmd1_scatter_groups_sva;
  reg while_case_28_lor_1_lpi_1_dfm;

  wire while_case_28_if_1_oelse_mux_1_nl;
  wire while_case_28_oelse_1_mux_1_nl;
  wire[31:0] while_case_28_if_1_oif_1_mul_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_ar_addr_rsc_dat_slave_process;
  assign nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_ar_addr_rsc_dat_slave_process
      = cmd1_ar_addr_sva;
  wire [31:0] nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_aw_addr_rsc_dat_slave_process;
  assign nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_aw_addr_rsc_dat_slave_process
      = cmd1_aw_addr_sva;
  wire [31:0] nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_total_len_rsc_dat_slave_process;
  assign nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_total_len_rsc_dat_slave_process
      = cmd1_total_len_sva;
  wire [31:0] nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_scatter_stride_rsc_dat_slave_process;
  assign nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_scatter_stride_rsc_dat_slave_process
      = cmd1_scatter_stride_sva;
  wire [15:0] nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_scatter_len_rsc_dat_slave_process;
  assign nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_scatter_len_rsc_dat_slave_process
      = cmd1_scatter_len_sva;
  wire [15:0] nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_scatter_groups_rsc_dat_slave_process;
  assign nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_scatter_groups_rsc_dat_slave_process
      = cmd1_scatter_groups_sva;
  wire [15:0] nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_dma_mode_rsc_dat_slave_process;
  assign nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_dma_mode_rsc_dat_slave_process
      = cmd1_dma_mode_sva;
  wire [1:0] nl_scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_inst_w_slave0_b_Push_mioi_idat_slave_process;
  assign nl_scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_inst_w_slave0_b_Push_mioi_idat_slave_process
      = {w_slave0_b_Push_mioi_idat_slave_process_1 , 1'b0};
  scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi scatter_gather_dma_slave_process_w_slave0_aw_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_slave0_aw_vld(w_slave0_aw_vld),
      .w_slave0_aw_rdy(w_slave0_aw_rdy),
      .w_slave0_aw_dat(w_slave0_aw_dat),
      .slave_process_wen(slave_process_wen),
      .w_slave0_aw_Pop_mioi_oswt(reg_w_slave0_w_Pop_mioi_iswt0_cse),
      .w_slave0_aw_Pop_mioi_wen_comp(w_slave0_aw_Pop_mioi_wen_comp),
      .w_slave0_aw_Pop_mioi_idat_mxwt(w_slave0_aw_Pop_mioi_idat_mxwt)
    );
  scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi scatter_gather_dma_slave_process_w_slave0_w_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_slave0_w_vld(w_slave0_w_vld),
      .w_slave0_w_rdy(w_slave0_w_rdy),
      .w_slave0_w_dat(w_slave0_w_dat),
      .slave_process_wen(slave_process_wen),
      .w_slave0_w_Pop_mioi_oswt(reg_w_slave0_w_Pop_mioi_iswt0_cse),
      .w_slave0_w_Pop_mioi_wen_comp(w_slave0_w_Pop_mioi_wen_comp),
      .w_slave0_w_Pop_mioi_idat_mxwt(w_slave0_w_Pop_mioi_idat_mxwt)
    );
  scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .dma_cmd_chan_vld(dma_cmd_chan_vld),
      .dma_cmd_chan_rdy(dma_cmd_chan_rdy),
      .dma_cmd_chan_dat(dma_cmd_chan_dat),
      .slave_process_wen(slave_process_wen),
      .dma_cmd_chan_Push_mioi_oswt(reg_dma_cmd_chan_Push_mioi_iswt0_cse),
      .dma_cmd_chan_Push_mioi_wen_comp(dma_cmd_chan_Push_mioi_wen_comp),
      .dma_cmd_chan_Push_mioi_m_ar_addr_rsc_dat_slave_process(nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_ar_addr_rsc_dat_slave_process[31:0]),
      .dma_cmd_chan_Push_mioi_m_aw_addr_rsc_dat_slave_process(nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_aw_addr_rsc_dat_slave_process[31:0]),
      .dma_cmd_chan_Push_mioi_m_total_len_rsc_dat_slave_process(nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_total_len_rsc_dat_slave_process[31:0]),
      .dma_cmd_chan_Push_mioi_m_scatter_stride_rsc_dat_slave_process(nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_scatter_stride_rsc_dat_slave_process[31:0]),
      .dma_cmd_chan_Push_mioi_m_scatter_len_rsc_dat_slave_process(nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_scatter_len_rsc_dat_slave_process[15:0]),
      .dma_cmd_chan_Push_mioi_m_scatter_groups_rsc_dat_slave_process(nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_scatter_groups_rsc_dat_slave_process[15:0]),
      .dma_cmd_chan_Push_mioi_m_dma_mode_rsc_dat_slave_process(nl_scatter_gather_dma_slave_process_dma_cmd_chan_Push_mioi_inst_dma_cmd_chan_Push_mioi_m_dma_mode_rsc_dat_slave_process[15:0]),
      .dma_cmd_chan_Push_mioi_oswt_pff(and_50_rmff)
    );
  scatter_gather_dma_slave_process_w_slave0_b_Push_mioi scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_slave0_b_vld(w_slave0_b_vld),
      .w_slave0_b_rdy(w_slave0_b_rdy),
      .w_slave0_b_dat(w_slave0_b_dat),
      .slave_process_wen(slave_process_wen),
      .w_slave0_b_Push_mioi_oswt(reg_w_slave0_b_Push_mioi_iswt0_cse),
      .w_slave0_b_Push_mioi_wen_comp(w_slave0_b_Push_mioi_wen_comp),
      .w_slave0_b_Push_mioi_idat_slave_process(nl_scatter_gather_dma_slave_process_w_slave0_b_Push_mioi_inst_w_slave0_b_Push_mioi_idat_slave_process[1:0])
    );
  scatter_gather_dma_slave_process_staller scatter_gather_dma_slave_process_staller_inst
      (
      .slave_process_wen(slave_process_wen),
      .w_slave0_aw_Pop_mioi_wen_comp(w_slave0_aw_Pop_mioi_wen_comp),
      .w_slave0_w_Pop_mioi_wen_comp(w_slave0_w_Pop_mioi_wen_comp),
      .dma_cmd_chan_Push_mioi_wen_comp(dma_cmd_chan_Push_mioi_wen_comp),
      .w_slave0_b_Push_mioi_wen_comp(w_slave0_b_Push_mioi_wen_comp)
    );
  scatter_gather_dma_slave_process_slave_process_fsm scatter_gather_dma_slave_process_slave_process_fsm_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .slave_process_wen(slave_process_wen),
      .fsm_output(fsm_output)
    );
  assign and_50_rmff = (~((while_case_28_if_1_oif_1_unequal_tmp | (cmd1_scatter_stride_sva[2:0]!=3'b000)
      | (cmd1_scatter_len_sva[2:0]!=3'b000)) & or_cse)) & (w_slave0_aw_Pop_mioi_idat_mxwt[29:0]==30'b000000000000000000000000011100)
      & (~((w_slave0_aw_Pop_mioi_idat_mxwt[31:30]!=2'b00) | while_case_28_if_while_case_28_if_or_1_tmp))
      & (fsm_output[1]);
  assign and_72_cse = while_switch_lp_nor_6_tmp & (w_slave0_aw_Pop_mioi_idat_mxwt[3:2]==2'b11);
  assign or_cse = (cmd1_dma_mode_sva!=16'b0000000000000000);
  assign while_case_28_if_while_case_28_if_or_1_tmp = (cmd1_total_len_sva[2:0]!=3'b000)
      | (cmd1_aw_addr_sva[2:0]!=3'b000) | (cmd1_ar_addr_sva[2:0]!=3'b000);
  assign while_case_28_if_1_lor_lpi_1_dfm_mx0w0 = (cmd1_scatter_stride_sva[2:0]!=3'b000)
      | (cmd1_scatter_len_sva[2:0]!=3'b000);
  assign while_case_28_if_1_oif_1_mul_nl = conv_u2u_32_32(cmd1_scatter_len_sva *
      cmd1_scatter_groups_sva);
  assign while_case_28_if_1_oif_1_unequal_tmp = while_case_28_if_1_oif_1_mul_nl !=
      cmd1_total_len_sva;
  assign while_switch_lp_while_switch_lp_nor_1_tmp = ~((w_slave0_aw_Pop_mioi_idat_mxwt!=32'b00000000000000000000000000000000));
  assign while_switch_lp_nor_1_tmp = ~((w_slave0_aw_Pop_mioi_idat_mxwt[31]) | (w_slave0_aw_Pop_mioi_idat_mxwt[30])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[29]) | (w_slave0_aw_Pop_mioi_idat_mxwt[28])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[27]) | (w_slave0_aw_Pop_mioi_idat_mxwt[26])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[25]) | (w_slave0_aw_Pop_mioi_idat_mxwt[24])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[23]) | (w_slave0_aw_Pop_mioi_idat_mxwt[22])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[21]) | (w_slave0_aw_Pop_mioi_idat_mxwt[20])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[19]) | (w_slave0_aw_Pop_mioi_idat_mxwt[18])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[17]) | (w_slave0_aw_Pop_mioi_idat_mxwt[16])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[15]) | (w_slave0_aw_Pop_mioi_idat_mxwt[14])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[13]) | (w_slave0_aw_Pop_mioi_idat_mxwt[12])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[11]) | (w_slave0_aw_Pop_mioi_idat_mxwt[10])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[9]) | (w_slave0_aw_Pop_mioi_idat_mxwt[8])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[7]) | (w_slave0_aw_Pop_mioi_idat_mxwt[6])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[5]) | (w_slave0_aw_Pop_mioi_idat_mxwt[4])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[3]) | (w_slave0_aw_Pop_mioi_idat_mxwt[1])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[0]));
  assign while_switch_lp_equal_tmp_7 = (w_slave0_aw_Pop_mioi_idat_mxwt[2]) & while_switch_lp_nor_1_tmp;
  assign while_switch_lp_nor_2_tmp = ~((w_slave0_aw_Pop_mioi_idat_mxwt[31]) | (w_slave0_aw_Pop_mioi_idat_mxwt[30])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[29]) | (w_slave0_aw_Pop_mioi_idat_mxwt[28])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[27]) | (w_slave0_aw_Pop_mioi_idat_mxwt[26])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[25]) | (w_slave0_aw_Pop_mioi_idat_mxwt[24])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[23]) | (w_slave0_aw_Pop_mioi_idat_mxwt[22])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[21]) | (w_slave0_aw_Pop_mioi_idat_mxwt[20])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[19]) | (w_slave0_aw_Pop_mioi_idat_mxwt[18])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[17]) | (w_slave0_aw_Pop_mioi_idat_mxwt[16])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[15]) | (w_slave0_aw_Pop_mioi_idat_mxwt[14])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[13]) | (w_slave0_aw_Pop_mioi_idat_mxwt[12])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[11]) | (w_slave0_aw_Pop_mioi_idat_mxwt[10])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[9]) | (w_slave0_aw_Pop_mioi_idat_mxwt[8])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[7]) | (w_slave0_aw_Pop_mioi_idat_mxwt[6])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[5]) | (w_slave0_aw_Pop_mioi_idat_mxwt[2])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[1]) | (w_slave0_aw_Pop_mioi_idat_mxwt[0]));
  assign while_switch_lp_equal_tmp_8 = (w_slave0_aw_Pop_mioi_idat_mxwt[4:3]==2'b11)
      & while_switch_lp_nor_2_tmp;
  assign while_switch_lp_nor_3_tmp = ~((w_slave0_aw_Pop_mioi_idat_mxwt[31]) | (w_slave0_aw_Pop_mioi_idat_mxwt[30])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[29]) | (w_slave0_aw_Pop_mioi_idat_mxwt[28])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[27]) | (w_slave0_aw_Pop_mioi_idat_mxwt[26])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[25]) | (w_slave0_aw_Pop_mioi_idat_mxwt[24])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[23]) | (w_slave0_aw_Pop_mioi_idat_mxwt[22])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[21]) | (w_slave0_aw_Pop_mioi_idat_mxwt[20])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[19]) | (w_slave0_aw_Pop_mioi_idat_mxwt[18])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[17]) | (w_slave0_aw_Pop_mioi_idat_mxwt[16])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[15]) | (w_slave0_aw_Pop_mioi_idat_mxwt[14])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[13]) | (w_slave0_aw_Pop_mioi_idat_mxwt[12])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[11]) | (w_slave0_aw_Pop_mioi_idat_mxwt[10])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[9]) | (w_slave0_aw_Pop_mioi_idat_mxwt[8])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[7]) | (w_slave0_aw_Pop_mioi_idat_mxwt[6])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[5]) | (w_slave0_aw_Pop_mioi_idat_mxwt[4])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[2]) | (w_slave0_aw_Pop_mioi_idat_mxwt[1])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[0]));
  assign while_switch_lp_equal_tmp_9 = (w_slave0_aw_Pop_mioi_idat_mxwt[3]) & while_switch_lp_nor_3_tmp;
  assign while_switch_lp_nor_4_tmp = ~((w_slave0_aw_Pop_mioi_idat_mxwt[31]) | (w_slave0_aw_Pop_mioi_idat_mxwt[30])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[29]) | (w_slave0_aw_Pop_mioi_idat_mxwt[28])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[27]) | (w_slave0_aw_Pop_mioi_idat_mxwt[26])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[25]) | (w_slave0_aw_Pop_mioi_idat_mxwt[24])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[23]) | (w_slave0_aw_Pop_mioi_idat_mxwt[22])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[21]) | (w_slave0_aw_Pop_mioi_idat_mxwt[20])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[19]) | (w_slave0_aw_Pop_mioi_idat_mxwt[18])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[17]) | (w_slave0_aw_Pop_mioi_idat_mxwt[16])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[15]) | (w_slave0_aw_Pop_mioi_idat_mxwt[14])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[13]) | (w_slave0_aw_Pop_mioi_idat_mxwt[12])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[11]) | (w_slave0_aw_Pop_mioi_idat_mxwt[10])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[9]) | (w_slave0_aw_Pop_mioi_idat_mxwt[8])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[7]) | (w_slave0_aw_Pop_mioi_idat_mxwt[6])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[5]) | (w_slave0_aw_Pop_mioi_idat_mxwt[3])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[2]) | (w_slave0_aw_Pop_mioi_idat_mxwt[1])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[0]));
  assign while_switch_lp_equal_tmp_10 = (w_slave0_aw_Pop_mioi_idat_mxwt[4]) & while_switch_lp_nor_4_tmp;
  assign while_switch_lp_nor_5_tmp = ~((w_slave0_aw_Pop_mioi_idat_mxwt[31]) | (w_slave0_aw_Pop_mioi_idat_mxwt[30])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[29]) | (w_slave0_aw_Pop_mioi_idat_mxwt[28])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[27]) | (w_slave0_aw_Pop_mioi_idat_mxwt[26])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[25]) | (w_slave0_aw_Pop_mioi_idat_mxwt[24])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[23]) | (w_slave0_aw_Pop_mioi_idat_mxwt[22])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[21]) | (w_slave0_aw_Pop_mioi_idat_mxwt[20])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[19]) | (w_slave0_aw_Pop_mioi_idat_mxwt[18])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[17]) | (w_slave0_aw_Pop_mioi_idat_mxwt[16])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[15]) | (w_slave0_aw_Pop_mioi_idat_mxwt[14])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[13]) | (w_slave0_aw_Pop_mioi_idat_mxwt[12])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[11]) | (w_slave0_aw_Pop_mioi_idat_mxwt[10])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[9]) | (w_slave0_aw_Pop_mioi_idat_mxwt[8])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[7]) | (w_slave0_aw_Pop_mioi_idat_mxwt[6])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[5]) | (w_slave0_aw_Pop_mioi_idat_mxwt[3])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[1]) | (w_slave0_aw_Pop_mioi_idat_mxwt[0]));
  assign while_switch_lp_equal_tmp_11 = (w_slave0_aw_Pop_mioi_idat_mxwt[4]) & (w_slave0_aw_Pop_mioi_idat_mxwt[2])
      & while_switch_lp_nor_5_tmp;
  assign while_switch_lp_nor_6_tmp = ~((w_slave0_aw_Pop_mioi_idat_mxwt[31]) | (w_slave0_aw_Pop_mioi_idat_mxwt[30])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[29]) | (w_slave0_aw_Pop_mioi_idat_mxwt[28])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[27]) | (w_slave0_aw_Pop_mioi_idat_mxwt[26])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[25]) | (w_slave0_aw_Pop_mioi_idat_mxwt[24])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[23]) | (w_slave0_aw_Pop_mioi_idat_mxwt[22])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[21]) | (w_slave0_aw_Pop_mioi_idat_mxwt[20])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[19]) | (w_slave0_aw_Pop_mioi_idat_mxwt[18])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[17]) | (w_slave0_aw_Pop_mioi_idat_mxwt[16])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[15]) | (w_slave0_aw_Pop_mioi_idat_mxwt[14])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[13]) | (w_slave0_aw_Pop_mioi_idat_mxwt[12])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[11]) | (w_slave0_aw_Pop_mioi_idat_mxwt[10])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[9]) | (w_slave0_aw_Pop_mioi_idat_mxwt[8])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[7]) | (w_slave0_aw_Pop_mioi_idat_mxwt[6])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[5]) | (w_slave0_aw_Pop_mioi_idat_mxwt[4])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[1]) | (w_slave0_aw_Pop_mioi_idat_mxwt[0]));
  assign or_dcpl_1 = (w_slave0_aw_Pop_mioi_idat_mxwt[31:30]!=2'b00);
  assign or_dcpl_5 = (w_slave0_aw_Pop_mioi_idat_mxwt[25:24]!=2'b00);
  assign or_dcpl_11 = (w_slave0_aw_Pop_mioi_idat_mxwt[19:18]!=2'b00);
  assign or_dcpl_17 = (w_slave0_aw_Pop_mioi_idat_mxwt[13:12]!=2'b00);
  assign or_dcpl_27 = ~((w_slave0_aw_Pop_mioi_idat_mxwt[3:2]==2'b11));
  assign or_dcpl_31 = or_dcpl_27 | (~ (w_slave0_aw_Pop_mioi_idat_mxwt[4])) | (w_slave0_aw_Pop_mioi_idat_mxwt[0])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[1]) | (w_slave0_aw_Pop_mioi_idat_mxwt[5])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[6]) | (w_slave0_aw_Pop_mioi_idat_mxwt[7])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[8]) | (w_slave0_aw_Pop_mioi_idat_mxwt[9])
      | (w_slave0_aw_Pop_mioi_idat_mxwt[10]) | (w_slave0_aw_Pop_mioi_idat_mxwt[11])
      | or_dcpl_17 | (w_slave0_aw_Pop_mioi_idat_mxwt[17:14]!=4'b0000) | or_dcpl_11
      | (w_slave0_aw_Pop_mioi_idat_mxwt[23:20]!=4'b0000) | or_dcpl_5 | (w_slave0_aw_Pop_mioi_idat_mxwt[29:26]!=4'b0000)
      | or_dcpl_1;
  assign and_dcpl_47 = (cmd1_dma_mode_sva==16'b0000000000000000);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_slave0_b_Push_mioi_idat_slave_process_1 <= 1'b0;
      reg_w_slave0_b_Push_mioi_iswt0_cse <= 1'b0;
      reg_dma_cmd_chan_Push_mioi_iswt0_cse <= 1'b0;
      reg_w_slave0_w_Pop_mioi_iswt0_cse <= 1'b0;
    end
    else if ( slave_process_wen ) begin
      w_slave0_b_Push_mioi_idat_slave_process_1 <= ((((while_case_28_if_1_oif_1_unequal_tmp
          | while_case_28_if_1_oelse_mux_1_nl) & or_cse) | while_case_28_oelse_1_mux_1_nl)
          & (~(while_switch_lp_while_switch_lp_nor_1_tmp | while_switch_lp_equal_tmp_7
          | while_switch_lp_equal_tmp_8 | while_switch_lp_equal_tmp_9 | while_switch_lp_equal_tmp_10
          | while_switch_lp_equal_tmp_11 | and_72_cse))) | (~(while_switch_lp_while_switch_lp_nor_1_tmp
          | while_switch_lp_equal_tmp_7 | while_switch_lp_equal_tmp_8 | while_switch_lp_equal_tmp_9
          | while_switch_lp_equal_tmp_10 | while_switch_lp_equal_tmp_11 | and_72_cse
          | ((w_slave0_aw_Pop_mioi_idat_mxwt==32'b00000000000000000000000000011100))));
      reg_w_slave0_b_Push_mioi_iswt0_cse <= fsm_output[1];
      reg_dma_cmd_chan_Push_mioi_iswt0_cse <= and_50_rmff;
      reg_w_slave0_w_Pop_mioi_iswt0_cse <= ~ (fsm_output[1]);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_case_28_lor_1_lpi_1_dfm <= 1'b0;
    end
    else if ( slave_process_wen & (~(or_dcpl_31 | (~ (fsm_output[1])))) ) begin
      while_case_28_lor_1_lpi_1_dfm <= while_case_28_if_while_case_28_if_or_1_tmp;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      cmd1_dma_mode_sva <= 16'b0000000000000000;
    end
    else if ( slave_process_wen & (w_slave0_aw_Pop_mioi_idat_mxwt[3]) & while_switch_lp_nor_2_tmp
        & (w_slave0_aw_Pop_mioi_idat_mxwt[4]) & (fsm_output[1]) ) begin
      cmd1_dma_mode_sva <= w_slave0_w_Pop_mioi_idat_mxwt[15:0];
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      cmd1_scatter_groups_sva <= 16'b0000000000000000;
    end
    else if ( slave_process_wen & (w_slave0_aw_Pop_mioi_idat_mxwt[2]) & while_switch_lp_nor_5_tmp
        & (w_slave0_aw_Pop_mioi_idat_mxwt[4]) & (fsm_output[1]) ) begin
      cmd1_scatter_groups_sva <= w_slave0_w_Pop_mioi_idat_mxwt[15:0];
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      cmd1_scatter_len_sva <= 16'b0000000000000000;
    end
    else if ( slave_process_wen & while_switch_lp_nor_4_tmp & (w_slave0_aw_Pop_mioi_idat_mxwt[4])
        & (fsm_output[1]) ) begin
      cmd1_scatter_len_sva <= w_slave0_w_Pop_mioi_idat_mxwt[15:0];
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      cmd1_scatter_stride_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( slave_process_wen & (~(or_dcpl_27 | (~ while_switch_lp_nor_6_tmp) |
        (~ (fsm_output[1])))) ) begin
      cmd1_scatter_stride_sva <= w_slave0_w_Pop_mioi_idat_mxwt;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      cmd1_total_len_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( slave_process_wen & (w_slave0_aw_Pop_mioi_idat_mxwt[3]) & while_switch_lp_nor_3_tmp
        & (fsm_output[1]) ) begin
      cmd1_total_len_sva <= w_slave0_w_Pop_mioi_idat_mxwt;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      cmd1_aw_addr_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( slave_process_wen & (w_slave0_aw_Pop_mioi_idat_mxwt[2]) & while_switch_lp_nor_1_tmp
        & (fsm_output[1]) ) begin
      cmd1_aw_addr_sva <= w_slave0_w_Pop_mioi_idat_mxwt;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      cmd1_ar_addr_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( slave_process_wen & while_switch_lp_while_switch_lp_nor_1_tmp & (fsm_output[1])
        ) begin
      cmd1_ar_addr_sva <= w_slave0_w_Pop_mioi_idat_mxwt;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_case_28_if_1_lor_lpi_1_dfm <= 1'b0;
    end
    else if ( slave_process_wen & (~(and_dcpl_47 | or_dcpl_27 | (~ (w_slave0_aw_Pop_mioi_idat_mxwt[4]))
        | (w_slave0_aw_Pop_mioi_idat_mxwt[0]) | (w_slave0_aw_Pop_mioi_idat_mxwt[1])
        | (w_slave0_aw_Pop_mioi_idat_mxwt[5]) | (w_slave0_aw_Pop_mioi_idat_mxwt[6])
        | (w_slave0_aw_Pop_mioi_idat_mxwt[7]) | (w_slave0_aw_Pop_mioi_idat_mxwt[8])
        | (w_slave0_aw_Pop_mioi_idat_mxwt[9]) | (w_slave0_aw_Pop_mioi_idat_mxwt[10])
        | (w_slave0_aw_Pop_mioi_idat_mxwt[11]) | or_dcpl_17 | (w_slave0_aw_Pop_mioi_idat_mxwt[17:14]!=4'b0000)
        | or_dcpl_11 | (w_slave0_aw_Pop_mioi_idat_mxwt[23:20]!=4'b0000) | or_dcpl_5
        | (w_slave0_aw_Pop_mioi_idat_mxwt[29:26]!=4'b0000) | or_dcpl_1 | while_case_28_if_while_case_28_if_or_1_tmp
        | (~ (fsm_output[1])))) ) begin
      while_case_28_if_1_lor_lpi_1_dfm <= while_case_28_if_1_lor_lpi_1_dfm_mx0w0;
    end
  end
  assign while_case_28_if_1_oelse_mux_1_nl = MUX_s_1_2_2(while_case_28_if_1_lor_lpi_1_dfm_mx0w0,
      while_case_28_if_1_lor_lpi_1_dfm, and_dcpl_47);
  assign while_case_28_oelse_1_mux_1_nl = MUX_s_1_2_2(while_case_28_if_while_case_28_if_or_1_tmp,
      while_case_28_lor_1_lpi_1_dfm, or_dcpl_31);

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_b_process
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_b_process (
  clk, rst_bar, b_in_vld, b_in_rdy, b_in_dat, b_chan_vld, b_chan_rdy, b_chan_dat,
      last_burst_chan_vld, last_burst_chan_rdy, last_burst_chan_dat
);
  input clk;
  input rst_bar;
  input b_in_vld;
  output b_in_rdy;
  input [5:0] b_in_dat;
  output b_chan_vld;
  input b_chan_rdy;
  output [5:0] b_chan_dat;
  input last_burst_chan_vld;
  output last_burst_chan_rdy;
  input last_burst_chan_dat;


  // Interconnect Declarations
  wire b_process_wen;
  wire b_process_wten;
  wire b_in_Pop_mioi_bawt;
  reg b_in_Pop_mioi_iswt0;
  wire b_in_Pop_mioi_wen_comp;
  wire [5:0] b_in_Pop_mioi_idat_mxwt;
  wire last_burst_chan_Pop_mioi_bawt;
  wire last_burst_chan_Pop_mioi_wen_comp;
  wire last_burst_chan_Pop_mioi_return_rsc_z_mxwt;
  wire b_chan_Push_mioi_bawt;
  reg b_chan_Push_mioi_iswt0;
  wire b_chan_Push_mioi_wen_comp;
  reg [1:0] b_chan_Push_mioi_idat_5_4;
  reg [3:0] b_chan_Push_mioi_idat_3_0;
  wire [1:0] fsm_output;
  wire and_dcpl;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire or_dcpl_3;
  wire or_dcpl_4;
  wire and_dcpl_10;
  wire and_dcpl_13;
  wire or_dcpl_10;
  wire or_tmp_6;
  wire while_stage_en_1_mx0w1;
  wire while_while_or_2_cse_1;
  wire while_while_or_1_cse_1;
  reg while_stage_v_1;
  reg while_stage_v_2;
  reg while_while_asn_mdf_sva_st_1;
  reg [3:0] comb_id_sva;
  reg id_valid_sva;
  wire while_while_and_1_tmp;
  wire while_while_if_1_and_cse;
  reg reg_last_burst_chan_Pop_mioi_iswt0_cse;
  wire while_and_cse;
  wire while_while_nand_cse;
  reg [1:0] comb_resp_sva;
  wire id_valid_sva_mx1;
  wire while_stage_v_2_mx0c1;
  wire [1:0] comb_resp_sva_mx0w0;

  wire[1:0] while_while_or_nl;
  wire[1:0] while_while_while_while_mux1h_nl;
  wire while_while_while_while_nor_nl;
  wire while_while_and_3_nl;
  wire mux_9_nl;
  wire while_while_not_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_inst_b_chan_Push_mioi_oswt_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_inst_b_chan_Push_mioi_oswt_unreg
      = b_chan_Push_mioi_bawt & while_while_asn_mdf_sva_st_1 & while_stage_v_2;
  wire [5:0] nl_axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_inst_b_chan_Push_mioi_idat;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_inst_b_chan_Push_mioi_idat
      = {b_chan_Push_mioi_idat_5_4 , b_chan_Push_mioi_idat_3_0};
  wire  nl_axi_axi4_segment_axi_cfg_standard_w_segment_b_process_staller_2_inst_b_process_flen_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_b_process_staller_2_inst_b_process_flen_unreg
      = ~(while_while_nand_cse | (while_stage_en_1_mx0w1 & (fsm_output[1])) | (while_stage_v_1
      & (~(while_stage_v_2 & and_dcpl)) & while_while_or_2_cse_1 & while_while_or_1_cse_1
      & (fsm_output[1])) | (while_stage_v_2 & while_while_or_1_cse_1 & (fsm_output[1])));
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_in_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .b_in_vld(b_in_vld),
      .b_in_rdy(b_in_rdy),
      .b_in_dat(b_in_dat),
      .b_in_Pop_mioi_oswt_unreg(or_tmp_6),
      .b_process_wen(b_process_wen),
      .b_process_wten(b_process_wten),
      .b_in_Pop_mioi_bawt(b_in_Pop_mioi_bawt),
      .b_in_Pop_mioi_iswt0(b_in_Pop_mioi_iswt0),
      .b_in_Pop_mioi_wen_comp(b_in_Pop_mioi_wen_comp),
      .b_in_Pop_mioi_idat_mxwt(b_in_Pop_mioi_idat_mxwt)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi
      axi_axi4_segment_axi_cfg_standard_w_segment_b_process_last_burst_chan_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_burst_chan_vld(last_burst_chan_vld),
      .last_burst_chan_rdy(last_burst_chan_rdy),
      .last_burst_chan_dat(last_burst_chan_dat),
      .last_burst_chan_Pop_mioi_oswt_unreg(and_dcpl_10),
      .b_process_wen(b_process_wen),
      .b_process_wten(b_process_wten),
      .last_burst_chan_Pop_mioi_bawt(last_burst_chan_Pop_mioi_bawt),
      .last_burst_chan_Pop_mioi_iswt0(reg_last_burst_chan_Pop_mioi_iswt0_cse),
      .last_burst_chan_Pop_mioi_wen_comp(last_burst_chan_Pop_mioi_wen_comp),
      .last_burst_chan_Pop_mioi_return_rsc_z_mxwt(last_burst_chan_Pop_mioi_return_rsc_z_mxwt),
      .last_burst_chan_Pop_mioi_iswt0_pff(or_tmp_6)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .b_chan_vld(b_chan_vld),
      .b_chan_rdy(b_chan_rdy),
      .b_chan_dat(b_chan_dat),
      .b_chan_Push_mioi_oswt_unreg(nl_axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_inst_b_chan_Push_mioi_oswt_unreg),
      .b_process_wen(b_process_wen),
      .b_process_wten(b_process_wten),
      .b_chan_Push_mioi_bawt(b_chan_Push_mioi_bawt),
      .b_chan_Push_mioi_iswt0(b_chan_Push_mioi_iswt0),
      .b_chan_Push_mioi_wen_comp(b_chan_Push_mioi_wen_comp),
      .b_chan_Push_mioi_idat(nl_axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_chan_Push_mioi_inst_b_chan_Push_mioi_idat[5:0])
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_staller_2 axi_axi4_segment_axi_cfg_standard_w_segment_b_process_staller_2_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .b_process_flen_unreg(nl_axi_axi4_segment_axi_cfg_standard_w_segment_b_process_staller_2_inst_b_process_flen_unreg),
      .b_process_wen(b_process_wen),
      .b_process_wten(b_process_wten),
      .b_in_Pop_mioi_wen_comp(b_in_Pop_mioi_wen_comp),
      .last_burst_chan_Pop_mioi_wen_comp(last_burst_chan_Pop_mioi_wen_comp),
      .b_chan_Push_mioi_wen_comp(b_chan_Push_mioi_wen_comp)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_process_fsm axi_axi4_segment_axi_cfg_standard_w_segment_b_process_b_process_fsm_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .b_process_wen(b_process_wen),
      .fsm_output(fsm_output)
    );
  assign while_while_nand_cse = ~((~ while_stage_en_1_mx0w1) & (fsm_output[1]));
  assign while_while_if_1_and_cse = b_process_wen & (~ and_dcpl_1) & last_burst_chan_Pop_mioi_bawt
      & last_burst_chan_Pop_mioi_return_rsc_z_mxwt & while_stage_v_1;
  assign while_and_cse = b_process_wen & (or_tmp_6 | and_dcpl_13);
  assign while_stage_en_1_mx0w1 = b_in_Pop_mioi_bawt & while_while_or_2_cse_1 & while_while_or_1_cse_1;
  assign id_valid_sva_mx1 = MUX_s_1_2_2(id_valid_sva, (~ last_burst_chan_Pop_mioi_return_rsc_z_mxwt),
      while_stage_v_1);
  assign while_while_not_nl = ~ last_burst_chan_Pop_mioi_return_rsc_z_mxwt;
  assign comb_resp_sva_mx0w0 = MUX_v_2_2_2(2'b00, comb_resp_sva, while_while_not_nl);
  assign while_while_or_2_cse_1 = last_burst_chan_Pop_mioi_bawt | (~ while_stage_v_1);
  assign while_while_or_1_cse_1 = b_chan_Push_mioi_bawt | (~(while_while_asn_mdf_sva_st_1
      & while_stage_v_2));
  assign and_dcpl = (~ b_chan_Push_mioi_bawt) & while_while_asn_mdf_sva_st_1;
  assign and_dcpl_1 = and_dcpl & while_stage_v_2;
  assign and_dcpl_2 = last_burst_chan_Pop_mioi_bawt & last_burst_chan_Pop_mioi_return_rsc_z_mxwt;
  assign or_dcpl_3 = b_chan_Push_mioi_bawt | (~ while_while_asn_mdf_sva_st_1);
  assign or_dcpl_4 = or_dcpl_3 | (~ while_stage_v_2);
  assign and_dcpl_10 = or_dcpl_4 & last_burst_chan_Pop_mioi_bawt & while_stage_v_1;
  assign and_dcpl_13 = or_dcpl_4 & last_burst_chan_Pop_mioi_bawt & (~ b_in_Pop_mioi_bawt)
      & while_stage_v_1;
  assign or_dcpl_10 = ~(last_burst_chan_Pop_mioi_bawt & while_stage_v_1);
  assign or_tmp_6 = or_dcpl_4 & b_in_Pop_mioi_bawt & while_while_or_2_cse_1 & (fsm_output[1]);
  assign while_stage_v_2_mx0c1 = or_dcpl_3 & while_stage_v_2 & or_dcpl_10;
  assign while_while_and_1_tmp = (comb_id_sva != (b_in_Pop_mioi_idat_mxwt[3:0]))
      & id_valid_sva_mx1;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      b_in_Pop_mioi_iswt0 <= 1'b0;
      b_chan_Push_mioi_iswt0 <= 1'b0;
      reg_last_burst_chan_Pop_mioi_iswt0_cse <= 1'b0;
    end
    else if ( b_process_wen ) begin
      b_in_Pop_mioi_iswt0 <= while_while_nand_cse;
      b_chan_Push_mioi_iswt0 <= or_dcpl_4 & and_dcpl_2 & while_stage_v_1;
      reg_last_burst_chan_Pop_mioi_iswt0_cse <= or_tmp_6;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      b_chan_Push_mioi_idat_3_0 <= 4'b0000;
      b_chan_Push_mioi_idat_5_4 <= 2'b00;
    end
    else if ( while_while_if_1_and_cse ) begin
      b_chan_Push_mioi_idat_3_0 <= comb_id_sva;
      b_chan_Push_mioi_idat_5_4 <= comb_resp_sva;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      id_valid_sva <= 1'b0;
    end
    else if ( b_process_wen & (~ (fsm_output[0])) ) begin
      id_valid_sva <= id_valid_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_stage_v_1 <= 1'b0;
      comb_resp_sva <= 2'b00;
    end
    else if ( while_and_cse ) begin
      while_stage_v_1 <= ~ and_dcpl_13;
      comb_resp_sva <= MUX_v_2_2_2(comb_resp_sva_mx0w0, while_while_or_nl, or_tmp_6);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_stage_v_2 <= 1'b0;
    end
    else if ( b_process_wen & (and_dcpl_10 | while_stage_v_2_mx0c1) ) begin
      while_stage_v_2 <= ~ while_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_while_asn_mdf_sva_st_1 <= 1'b0;
    end
    else if ( b_process_wen & (~(and_dcpl_1 | or_dcpl_10)) ) begin
      while_while_asn_mdf_sva_st_1 <= last_burst_chan_Pop_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      comb_id_sva <= 4'b0000;
    end
    else if ( b_process_wen & (~(mux_9_nl | and_dcpl_1 | (~ b_in_Pop_mioi_bawt)))
        ) begin
      comb_id_sva <= b_in_Pop_mioi_idat_mxwt[3:0];
    end
  end
  assign while_while_while_while_nor_nl = ~(while_stage_v_1 | while_while_and_1_tmp);
  assign while_while_and_3_nl = while_stage_v_1 & (~ while_while_and_1_tmp);
  assign while_while_while_while_mux1h_nl = MUX1HOT_v_2_3_2(comb_resp_sva, comb_resp_sva_mx0w0,
      2'b10, {while_while_while_while_nor_nl , while_while_and_3_nl , while_while_and_1_tmp});
  assign while_while_or_nl = while_while_while_while_mux1h_nl | (b_in_Pop_mioi_idat_mxwt[5:4]);
  assign mux_9_nl = MUX_s_1_2_2(id_valid_sva, (~ and_dcpl_2), while_stage_v_1);

  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_w_process
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_w_process (
  clk, rst_bar, w_out_vld, w_out_rdy, w_out_dat, w_chan_vld, w_chan_rdy, w_chan_dat,
      last_bit_chan_vld, last_bit_chan_rdy, last_bit_chan_dat
);
  input clk;
  input rst_bar;
  output w_out_vld;
  input w_out_rdy;
  output [72:0] w_out_dat;
  input w_chan_vld;
  output w_chan_rdy;
  input [72:0] w_chan_dat;
  input last_bit_chan_vld;
  output last_bit_chan_rdy;
  input last_bit_chan_dat;


  // Interconnect Declarations
  wire w_process_wen;
  wire w_process_wten;
  wire w_chan_Pop_mioi_bawt;
  reg w_chan_Pop_mioi_iswt0;
  wire w_chan_Pop_mioi_wen_comp;
  wire [71:0] w_chan_Pop_mioi_idat_mxwt;
  wire last_bit_chan_Pop_mioi_bawt;
  wire last_bit_chan_Pop_mioi_wen_comp;
  wire last_bit_chan_Pop_mioi_return_rsc_z_mxwt;
  wire w_out_Push_mioi_bawt;
  wire w_out_Push_mioi_wen_comp;
  reg [7:0] w_out_Push_mioi_idat_72_65;
  reg w_out_Push_mioi_idat_64;
  reg [63:0] w_out_Push_mioi_idat_63_0;
  wire [1:0] fsm_output;
  wire or_dcpl;
  wire and_dcpl;
  wire and_dcpl_2;
  wire and_dcpl_5;
  wire or_tmp_4;
  wire while_stage_en_1_mx0w1;
  wire while_while_or_1_cse_1;
  wire while_while_or_cse_1;
  reg while_stage_v_1;
  reg while_stage_v_2;
  wire while_and_cse;
  reg reg_w_out_Push_mioi_iswt0_cse;
  reg reg_last_bit_chan_Pop_mioi_iswt0_cse;
  wire while_nand_cse;
  reg [7:0] while_slc_assocmrg_72_65_itm_1;
  reg [63:0] while_slc_assocmrg_63_0_itm_1;
  wire while_stage_v_1_mx0c1;
  wire while_stage_v_2_mx0c1;
  wire while_and_11_cse;


  // Interconnect Declarations for Component Instantiations 
  wire [72:0] nl_axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_inst_w_out_Push_mioi_idat;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_inst_w_out_Push_mioi_idat
      = {w_out_Push_mioi_idat_72_65 , w_out_Push_mioi_idat_64 , w_out_Push_mioi_idat_63_0};
  wire  nl_axi_axi4_segment_axi_cfg_standard_w_segment_w_process_staller_1_inst_w_process_flen_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_w_process_staller_1_inst_w_process_flen_unreg
      = ~(while_nand_cse | (while_stage_en_1_mx0w1 & (fsm_output[1])) | (while_stage_v_1
      & (~(while_stage_v_2 & (~ w_out_Push_mioi_bawt))) & while_while_or_1_cse_1
      & while_while_or_cse_1 & (fsm_output[1])) | (while_stage_v_2 & while_while_or_cse_1
      & (fsm_output[1])));
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_chan_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_chan_vld(w_chan_vld),
      .w_chan_rdy(w_chan_rdy),
      .w_chan_dat(w_chan_dat),
      .w_chan_Pop_mioi_oswt_unreg(or_tmp_4),
      .w_process_wen(w_process_wen),
      .w_process_wten(w_process_wten),
      .w_chan_Pop_mioi_bawt(w_chan_Pop_mioi_bawt),
      .w_chan_Pop_mioi_iswt0(w_chan_Pop_mioi_iswt0),
      .w_chan_Pop_mioi_wen_comp(w_chan_Pop_mioi_wen_comp),
      .w_chan_Pop_mioi_idat_mxwt(w_chan_Pop_mioi_idat_mxwt)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi axi_axi4_segment_axi_cfg_standard_w_segment_w_process_last_bit_chan_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_bit_chan_vld(last_bit_chan_vld),
      .last_bit_chan_rdy(last_bit_chan_rdy),
      .last_bit_chan_dat(last_bit_chan_dat),
      .last_bit_chan_Pop_mioi_oswt_unreg(and_dcpl_2),
      .w_process_wen(w_process_wen),
      .w_process_wten(w_process_wten),
      .last_bit_chan_Pop_mioi_bawt(last_bit_chan_Pop_mioi_bawt),
      .last_bit_chan_Pop_mioi_iswt0(reg_last_bit_chan_Pop_mioi_iswt0_cse),
      .last_bit_chan_Pop_mioi_wen_comp(last_bit_chan_Pop_mioi_wen_comp),
      .last_bit_chan_Pop_mioi_return_rsc_z_mxwt(last_bit_chan_Pop_mioi_return_rsc_z_mxwt),
      .last_bit_chan_Pop_mioi_iswt0_pff(or_tmp_4)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_out_vld(w_out_vld),
      .w_out_rdy(w_out_rdy),
      .w_out_dat(w_out_dat),
      .w_out_Push_mioi_oswt_unreg(and_dcpl_5),
      .w_process_wen(w_process_wen),
      .w_process_wten(w_process_wten),
      .w_out_Push_mioi_bawt(w_out_Push_mioi_bawt),
      .w_out_Push_mioi_iswt0(reg_w_out_Push_mioi_iswt0_cse),
      .w_out_Push_mioi_wen_comp(w_out_Push_mioi_wen_comp),
      .w_out_Push_mioi_idat(nl_axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_out_Push_mioi_inst_w_out_Push_mioi_idat[72:0])
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_staller_1 axi_axi4_segment_axi_cfg_standard_w_segment_w_process_staller_1_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_process_flen_unreg(nl_axi_axi4_segment_axi_cfg_standard_w_segment_w_process_staller_1_inst_w_process_flen_unreg),
      .w_process_wen(w_process_wen),
      .w_process_wten(w_process_wten),
      .w_chan_Pop_mioi_wen_comp(w_chan_Pop_mioi_wen_comp),
      .last_bit_chan_Pop_mioi_wen_comp(last_bit_chan_Pop_mioi_wen_comp),
      .w_out_Push_mioi_wen_comp(w_out_Push_mioi_wen_comp)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_process_fsm axi_axi4_segment_axi_cfg_standard_w_segment_w_process_w_process_fsm_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_process_wen(w_process_wen),
      .fsm_output(fsm_output)
    );
  assign while_nand_cse = ~((~ while_stage_en_1_mx0w1) & (fsm_output[1]));
  assign while_and_cse = w_process_wen & (~(and_dcpl | or_dcpl));
  assign while_and_11_cse = w_process_wen & (~(and_dcpl | ((~ last_bit_chan_Pop_mioi_bawt)
      & while_stage_v_1)));
  assign while_stage_en_1_mx0w1 = w_chan_Pop_mioi_bawt & while_while_or_1_cse_1 &
      while_while_or_cse_1;
  assign while_while_or_1_cse_1 = last_bit_chan_Pop_mioi_bawt | (~ while_stage_v_1);
  assign while_while_or_cse_1 = w_out_Push_mioi_bawt | (~ while_stage_v_2);
  assign or_dcpl = ~(last_bit_chan_Pop_mioi_bawt & while_stage_v_1);
  assign and_dcpl = (~ w_out_Push_mioi_bawt) & while_stage_v_2;
  assign and_dcpl_2 = while_while_or_cse_1 & while_stage_v_1 & last_bit_chan_Pop_mioi_bawt;
  assign and_dcpl_5 = w_out_Push_mioi_bawt & while_stage_v_2;
  assign or_tmp_4 = while_while_or_cse_1 & while_while_or_1_cse_1 & w_chan_Pop_mioi_bawt
      & (fsm_output[1]);
  assign while_stage_v_1_mx0c1 = while_while_or_cse_1 & last_bit_chan_Pop_mioi_bawt
      & while_stage_v_1 & (~ w_chan_Pop_mioi_bawt);
  assign while_stage_v_2_mx0c1 = and_dcpl_5 & or_dcpl;
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_chan_Pop_mioi_iswt0 <= 1'b0;
      reg_w_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_last_bit_chan_Pop_mioi_iswt0_cse <= 1'b0;
    end
    else if ( w_process_wen ) begin
      w_chan_Pop_mioi_iswt0 <= while_nand_cse;
      reg_w_out_Push_mioi_iswt0_cse <= and_dcpl_2;
      reg_last_bit_chan_Pop_mioi_iswt0_cse <= or_tmp_4;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      w_out_Push_mioi_idat_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      w_out_Push_mioi_idat_64 <= 1'b0;
      w_out_Push_mioi_idat_72_65 <= 8'b00000000;
    end
    else if ( while_and_cse ) begin
      w_out_Push_mioi_idat_63_0 <= while_slc_assocmrg_63_0_itm_1;
      w_out_Push_mioi_idat_64 <= last_bit_chan_Pop_mioi_return_rsc_z_mxwt;
      w_out_Push_mioi_idat_72_65 <= while_slc_assocmrg_72_65_itm_1;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_stage_v_1 <= 1'b0;
    end
    else if ( w_process_wen & (or_tmp_4 | while_stage_v_1_mx0c1) ) begin
      while_stage_v_1 <= ~ while_stage_v_1_mx0c1;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_slc_assocmrg_72_65_itm_1 <= 8'b00000000;
      while_slc_assocmrg_63_0_itm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( while_and_11_cse ) begin
      while_slc_assocmrg_72_65_itm_1 <= w_chan_Pop_mioi_idat_mxwt[71:64];
      while_slc_assocmrg_63_0_itm_1 <= w_chan_Pop_mioi_idat_mxwt[63:0];
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_stage_v_2 <= 1'b0;
    end
    else if ( w_process_wen & (and_dcpl_2 | while_stage_v_2_mx0c1) ) begin
      while_stage_v_2 <= ~ while_stage_v_2_mx0c1;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process (
  clk, rst_bar, aw_out_vld, aw_out_rdy, aw_out_dat, ex_aw_chan_vld, ex_aw_chan_rdy,
      ex_aw_chan_dat, last_bit_chan_vld, last_bit_chan_rdy, last_bit_chan_dat, last_burst_chan_vld,
      last_burst_chan_rdy, last_burst_chan_dat
);
  input clk;
  input rst_bar;
  output aw_out_vld;
  input aw_out_rdy;
  output [43:0] aw_out_dat;
  input ex_aw_chan_vld;
  output ex_aw_chan_rdy;
  input [75:0] ex_aw_chan_dat;
  output last_bit_chan_vld;
  input last_bit_chan_rdy;
  output last_bit_chan_dat;
  output last_burst_chan_vld;
  input last_burst_chan_rdy;
  output last_burst_chan_dat;


  // Interconnect Declarations
  wire ex_aw_process_wen;
  wire ex_aw_process_wten;
  wire ex_aw_chan_Pop_mioi_bawt;
  reg ex_aw_chan_Pop_mioi_iswt0;
  wire ex_aw_chan_Pop_mioi_wen_comp;
  wire [67:0] ex_aw_chan_Pop_mioi_idat_mxwt;
  wire aw_out_Push_mioi_bawt;
  reg aw_out_Push_mioi_iswt0;
  wire aw_out_Push_mioi_wen_comp;
  wire last_bit_chan_Push_mioi_bawt;
  reg last_bit_chan_Push_mioi_iswt0;
  wire last_bit_chan_Push_mioi_wen_comp;
  reg last_bit_chan_Push_mioi_m_rsc_dat;
  wire last_burst_chan_Push_mioi_bawt;
  reg last_burst_chan_Push_mioi_iswt0;
  wire last_burst_chan_Push_mioi_wen_comp;
  reg last_burst_chan_Push_mioi_m_rsc_dat;
  reg [6:0] aw_out_Push_mioi_idat_6_0;
  reg [24:0] aw_out_Push_mioi_idat_35_11;
  reg [3:0] aw_out_Push_mioi_idat_10_7;
  reg [4:0] aw_out_Push_mioi_idat_40_36;
  wire [1:0] fsm_output;
  wire [4:0] while_while_if_1_mux_2_tmp;
  wire [9:0] operator_8_false_1_acc_tmp;
  wire [10:0] nl_operator_8_false_1_acc_tmp;
  wire while_while_while_while_or_tmp;
  wire or_dcpl_4;
  wire nand_tmp_6;
  wire and_dcpl_4;
  wire and_dcpl_7;
  wire or_dcpl_21;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_18;
  wire and_dcpl_19;
  wire and_dcpl_22;
  wire and_dcpl_24;
  wire and_dcpl_37;
  wire or_tmp_78;
  wire while_stage_en_1_mx0w1;
  wire while_while_last_burst_lpi_1_dfm_2_mx0;
  wire while_while_while_last_sva_mx1w0;
  wire [7:0] while_while_aw_len_lpi_1_dfm_3_mx0;
  reg while_while_asn_itm;
  wire while_or_cse_1;
  wire while_or_1_cse_1;
  wire while_or_2_cse_1;
  reg while_stage_v_1;
  reg while_while_while_last_sva_st_1;
  reg exitL_exit_while_while_while_lpi_1_dfm_st_1;
  reg exitL_exit_while_while_sva;
  reg [7:0] while_while_aw_len_lpi_1;
  reg while_while_last_burst_lpi_1_dfm_2;
  reg exit_while_while_lpi_1_dfm_1;
  reg exitL_exit_while_while_while_lpi_1;
  wire or_56_cse;
  wire while_while_and_1_cse;
  wire or_49_cse;
  wire while_while_and_cse;
  wire or_132_cse;
  wire or_19_cse;
  wire nand_16_cse;
  wire or_106_cse;
  wire or_5_cse;
  wire [7:0] while_while_aw_len_sva_4;
  wire [8:0] nl_while_while_aw_len_sva_4;
  wire mux_30_cse;
  wire and_136_cse;
  wire while_ex_addr_and_4_cse;
  wire and_137_cse;
  wire while_while_aw_out_write_reset_check_ResetChecker_nand_cse;
  wire and_15_cse;
  wire nand_1_cse;
  wire while_while_while_mux_rmff;
  wire while_while_mux_5_rmff;
  wire and_103_rmff;
  wire or_tmp_92;
  wire [28:0] z_out;
  reg [24:0] while_ex_addr_31_3_lpi_1_28_4;
  reg [3:0] while_ex_addr_31_3_lpi_1_3_0;
  reg [27:0] while_ex_ex_len_lpi_1_31_4;
  reg [3:0] while_ex_ex_len_lpi_1_3_0;
  reg [6:0] assocmrg_lpi_1_dfm_6_0;
  wire while_while_if_1_if_while_while_if_1_if_nor_mx1w0;
  wire exit_while_while_lpi_1_dfm_1_mx0w0;
  wire while_stage_v_1_mx0c1;
  wire [4:0] while_while_aw_len_sva_2_4_0_2;
  wire [5:0] nl_while_while_aw_len_sva_2_4_0_2;
  wire [3:0] while_while_while_while_or_3_psp_1;
  wire [4:0] while_while_if_1_mux_2_psp_mx0;
  wire [24:0] while_ex_addr_31_3_lpi_1_dfm_28_4_mx0;
  wire [3:0] while_ex_addr_31_3_lpi_1_dfm_3_0_mx0;
  wire [3:0] while_ex_ex_len_lpi_1_dfm_3_0_mx0;
  wire [27:0] while_ex_ex_len_lpi_1_dfm_31_4_mx0;
  wire [28:0] while_ex_addr_31_3_sva_5;
  wire [29:0] nl_while_ex_addr_31_3_sva_5;
  wire [31:0] while_ex_ex_len_sva_4;
  wire [32:0] nl_while_ex_ex_len_sva_4;
  wire [27:0] while_ex_ex_len_lpi_1_dfm_1_31_4_1;
  wire [3:0] while_ex_ex_len_lpi_1_dfm_1_3_0_1;
  wire while_while_while_asn_12;
  wire and_28_rgt;
  wire and_78_rgt;
  wire while_while_and_9_cse;
  wire while_ex_addr_and_cse;
  wire operator_32_false_acc_itm_28_1;

  wire mux_29_nl;
  wire mux_28_nl;
  wire mux_27_nl;
  wire nor_10_nl;
  wire mux_26_nl;
  wire mux_25_nl;
  wire mux_24_nl;
  wire or_58_nl;
  wire and_18_nl;
  wire mux_23_nl;
  wire nand_5_nl;
  wire or_50_nl;
  wire nor_13_nl;
  wire nor_14_nl;
  wire while_while_if_1_if_mux1h_nl;
  wire and_41_nl;
  wire and_44_nl;
  wire and_48_nl;
  wire or_85_nl;
  wire mux_32_nl;
  wire mux_31_nl;
  wire or_84_nl;
  wire or_83_nl;
  wire or_81_nl;
  wire mux_34_nl;
  wire nor_9_nl;
  wire while_while_while_last_mux_nl;
  wire and_74_nl;
  wire and_75_nl;
  wire[28:0] operator_32_false_acc_nl;
  wire[29:0] nl_operator_32_false_acc_nl;
  wire while_while_aw_len_and_nl;
  wire while_while_aw_len_and_1_nl;
  wire nand_25_nl;
  wire[24:0] while_while_mux_13_nl;
  wire[3:0] while_while_mux_12_nl;
  wire[27:0] operator_32_false_acc_nl_1;
  wire[28:0] nl_operator_32_false_acc_nl_1;
  wire while_while_not_26_nl;
  wire while_while_not_22_nl;
  wire[29:0] acc_nl;
  wire[30:0] nl_acc_nl;
  wire[28:0] operator_8_false_mux_2_nl;
  wire operator_8_false_operator_8_false_nand_1_nl;
  wire[3:0] operator_8_false_mux_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_inst_ex_aw_chan_Pop_mioi_oswt_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_inst_ex_aw_chan_Pop_mioi_oswt_unreg
      = while_while_aw_out_write_reset_check_ResetChecker_nand_cse & while_while_asn_itm
      & ex_aw_chan_Pop_mioi_bawt & (fsm_output[1]);
  wire  nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_inst_aw_out_Push_mioi_oswt_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_inst_aw_out_Push_mioi_oswt_unreg
      = or_132_cse & aw_out_Push_mioi_bawt & last_bit_chan_Push_mioi_bawt & exitL_exit_while_while_while_lpi_1_dfm_st_1
      & while_stage_v_1;
  wire [43:0] nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_inst_aw_out_Push_mioi_idat;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_inst_aw_out_Push_mioi_idat
      = signext_44_41({aw_out_Push_mioi_idat_40_36 , aw_out_Push_mioi_idat_35_11
      , aw_out_Push_mioi_idat_10_7 , aw_out_Push_mioi_idat_6_0});
  wire  nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_inst_last_bit_chan_Push_mioi_oswt_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_inst_last_bit_chan_Push_mioi_oswt_unreg
      = and_dcpl_37 & last_bit_chan_Push_mioi_bawt & while_stage_v_1;
  wire  nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_inst_last_burst_chan_Push_mioi_oswt_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_inst_last_burst_chan_Push_mioi_oswt_unreg
      = and_15_cse & last_burst_chan_Push_mioi_bawt & while_while_while_last_sva_st_1
      & while_stage_v_1;
  wire  nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_inst_last_burst_chan_Push_mioi_iswt0_pff;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_inst_last_burst_chan_Push_mioi_iswt0_pff
      = and_103_rmff;
  wire  nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_staller_inst_ex_aw_process_flen_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_staller_inst_ex_aw_process_flen_unreg
      = ~((~((~ while_stage_en_1_mx0w1) & (fsm_output[1]))) | (while_stage_en_1_mx0w1
      & (fsm_output[1])) | (while_stage_v_1 & while_or_cse_1 & while_or_1_cse_1 &
      while_or_2_cse_1 & (fsm_output[1])));
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_aw_chan_vld(ex_aw_chan_vld),
      .ex_aw_chan_rdy(ex_aw_chan_rdy),
      .ex_aw_chan_dat(ex_aw_chan_dat),
      .ex_aw_process_wen(ex_aw_process_wen),
      .ex_aw_process_wten(ex_aw_process_wten),
      .ex_aw_chan_Pop_mioi_oswt_unreg(nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_chan_Pop_mioi_inst_ex_aw_chan_Pop_mioi_oswt_unreg),
      .ex_aw_chan_Pop_mioi_bawt(ex_aw_chan_Pop_mioi_bawt),
      .ex_aw_chan_Pop_mioi_iswt0(ex_aw_chan_Pop_mioi_iswt0),
      .ex_aw_chan_Pop_mioi_wen_comp(ex_aw_chan_Pop_mioi_wen_comp),
      .ex_aw_chan_Pop_mioi_idat_mxwt(ex_aw_chan_Pop_mioi_idat_mxwt)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .aw_out_vld(aw_out_vld),
      .aw_out_rdy(aw_out_rdy),
      .aw_out_dat(aw_out_dat),
      .ex_aw_process_wen(ex_aw_process_wen),
      .ex_aw_process_wten(ex_aw_process_wten),
      .aw_out_Push_mioi_oswt_unreg(nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_inst_aw_out_Push_mioi_oswt_unreg),
      .aw_out_Push_mioi_bawt(aw_out_Push_mioi_bawt),
      .aw_out_Push_mioi_iswt0(aw_out_Push_mioi_iswt0),
      .aw_out_Push_mioi_wen_comp(aw_out_Push_mioi_wen_comp),
      .aw_out_Push_mioi_idat(nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_aw_out_Push_mioi_inst_aw_out_Push_mioi_idat[43:0])
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_bit_chan_vld(last_bit_chan_vld),
      .last_bit_chan_rdy(last_bit_chan_rdy),
      .last_bit_chan_dat(last_bit_chan_dat),
      .ex_aw_process_wen(ex_aw_process_wen),
      .ex_aw_process_wten(ex_aw_process_wten),
      .last_bit_chan_Push_mioi_oswt_unreg(nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_bit_chan_Push_mioi_inst_last_bit_chan_Push_mioi_oswt_unreg),
      .last_bit_chan_Push_mioi_bawt(last_bit_chan_Push_mioi_bawt),
      .last_bit_chan_Push_mioi_iswt0(last_bit_chan_Push_mioi_iswt0),
      .last_bit_chan_Push_mioi_wen_comp(last_bit_chan_Push_mioi_wen_comp),
      .last_bit_chan_Push_mioi_m_rsc_dat(while_while_while_mux_rmff),
      .last_bit_chan_Push_mioi_iswt0_pff(or_tmp_78)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi
      axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .last_burst_chan_vld(last_burst_chan_vld),
      .last_burst_chan_rdy(last_burst_chan_rdy),
      .last_burst_chan_dat(last_burst_chan_dat),
      .ex_aw_process_wen(ex_aw_process_wen),
      .ex_aw_process_wten(ex_aw_process_wten),
      .last_burst_chan_Push_mioi_oswt_unreg(nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_inst_last_burst_chan_Push_mioi_oswt_unreg),
      .last_burst_chan_Push_mioi_bawt(last_burst_chan_Push_mioi_bawt),
      .last_burst_chan_Push_mioi_iswt0(last_burst_chan_Push_mioi_iswt0),
      .last_burst_chan_Push_mioi_wen_comp(last_burst_chan_Push_mioi_wen_comp),
      .last_burst_chan_Push_mioi_m_rsc_dat(while_while_mux_5_rmff),
      .last_burst_chan_Push_mioi_iswt0_pff(nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_last_burst_chan_Push_mioi_inst_last_burst_chan_Push_mioi_iswt0_pff)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_staller axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_staller_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_aw_process_wen(ex_aw_process_wen),
      .ex_aw_process_wten(ex_aw_process_wten),
      .ex_aw_chan_Pop_mioi_wen_comp(ex_aw_chan_Pop_mioi_wen_comp),
      .aw_out_Push_mioi_wen_comp(aw_out_Push_mioi_wen_comp),
      .last_bit_chan_Push_mioi_wen_comp(last_bit_chan_Push_mioi_wen_comp),
      .last_burst_chan_Push_mioi_wen_comp(last_burst_chan_Push_mioi_wen_comp),
      .ex_aw_process_flen_unreg(nl_axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_staller_inst_ex_aw_process_flen_unreg)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_process_fsm axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_ex_aw_process_fsm_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_aw_process_wen(ex_aw_process_wen),
      .fsm_output(fsm_output)
    );
  assign or_56_cse = (operator_8_false_1_acc_tmp[3:0]!=4'b0000);
  assign or_49_cse = (~ while_while_asn_itm) | ex_aw_chan_Pop_mioi_bawt;
  assign while_while_and_cse = ex_aw_process_wen & (~(or_dcpl_21 | (fsm_output[0])));
  assign while_while_and_1_cse = ex_aw_process_wen & (~ (fsm_output[0]));
  assign and_137_cse = or_56_cse & (operator_8_false_1_acc_tmp[9]);
  assign and_28_rgt = (~(and_137_cse | and_dcpl_7)) & or_49_cse & or_5_cse;
  assign while_while_and_9_cse = while_while_and_1_cse & ((and_dcpl_15 & exitL_exit_while_while_sva)
      | and_dcpl_18);
  assign nand_16_cse = ~(last_bit_chan_Push_mioi_bawt & or_19_cse & or_132_cse);
  assign nor_13_nl = ~((while_while_aw_len_lpi_1!=8'b00000000));
  assign nor_14_nl = ~((while_while_aw_len_sva_4!=8'b00000000) | nand_16_cse);
  assign mux_30_cse = MUX_s_1_2_2(nor_13_nl, nor_14_nl, while_stage_v_1);
  assign and_136_cse = while_stage_v_1 & nand_16_cse;
  assign and_41_nl = and_dcpl_24 & and_dcpl_22 & and_dcpl_19 & (operator_8_false_1_acc_tmp[9]);
  assign and_44_nl = and_dcpl_24 & and_dcpl_22 & and_dcpl_19 & (~ (operator_8_false_1_acc_tmp[9]));
  assign and_48_nl = mux_30_cse & or_49_cse & and_dcpl_14;
  assign or_84_nl = (while_while_aw_len_lpi_1!=8'b00000000);
  assign or_83_nl = (while_while_aw_len_sva_4!=8'b00000000) | nand_16_cse;
  assign mux_31_nl = MUX_s_1_2_2(or_84_nl, or_83_nl, while_stage_v_1);
  assign or_81_nl = (while_while_if_1_mux_2_tmp!=5'b00000) | and_136_cse;
  assign mux_32_nl = MUX_s_1_2_2(mux_31_nl, or_81_nl, while_while_while_while_or_tmp);
  assign or_85_nl = mux_32_nl | and_dcpl_4;
  assign while_while_if_1_if_mux1h_nl = MUX1HOT_s_1_4_2(while_while_if_1_if_while_while_if_1_if_nor_mx1w0,
      (~ operator_32_false_acc_itm_28_1), while_while_last_burst_lpi_1_dfm_2, last_burst_chan_Push_mioi_m_rsc_dat,
      {and_41_nl , and_44_nl , and_48_nl , or_85_nl});
  assign while_while_mux_5_rmff = MUX_s_1_2_2(while_while_if_1_if_mux1h_nl, last_burst_chan_Push_mioi_m_rsc_dat,
      fsm_output[0]);
  assign nor_9_nl = ~((while_while_if_1_mux_2_tmp!=5'b00000) | and_136_cse);
  assign mux_34_nl = MUX_s_1_2_2(mux_30_cse, nor_9_nl, while_while_while_while_or_tmp);
  assign and_103_rmff = mux_34_nl & or_49_cse & (fsm_output[1]);
  assign while_while_while_last_mux_nl = MUX_s_1_2_2(while_while_while_last_sva_mx1w0,
      last_bit_chan_Push_mioi_m_rsc_dat, or_dcpl_21);
  assign while_while_while_mux_rmff = MUX_s_1_2_2(while_while_while_last_mux_nl,
      last_bit_chan_Push_mioi_m_rsc_dat, fsm_output[0]);
  assign or_132_cse = (~ while_while_while_last_sva_st_1) | last_burst_chan_Push_mioi_bawt;
  assign and_15_cse = last_bit_chan_Push_mioi_bawt & or_19_cse;
  assign nand_1_cse = ~(while_stage_v_1 & nand_16_cse);
  assign and_78_rgt = or_5_cse & or_49_cse;
  assign while_ex_addr_and_4_cse = while_while_while_asn_12 & (~ or_dcpl_21);
  assign while_ex_addr_and_cse = ex_aw_process_wen & (((~ and_137_cse) & while_while_while_while_or_tmp
      & (~ or_dcpl_21)) | while_ex_addr_and_4_cse);
  assign while_while_if_1_if_while_while_if_1_if_nor_mx1w0 = ~(operator_32_false_acc_itm_28_1
      | or_56_cse);
  assign while_while_while_last_sva_mx1w0 = ~((while_while_aw_len_lpi_1_dfm_3_mx0!=8'b00000000));
  assign or_106_cse = (~((~(exitL_exit_while_while_while_lpi_1_dfm_st_1 & (~ aw_out_Push_mioi_bawt)))
      & last_bit_chan_Push_mioi_bawt)) | ((~ last_burst_chan_Push_mioi_bawt) & while_while_while_last_sva_st_1);
  assign while_while_aw_out_write_reset_check_ResetChecker_nand_cse = ~(while_stage_v_1
      & or_106_cse);
  assign while_stage_en_1_mx0w1 = or_49_cse & while_or_cse_1 & while_or_1_cse_1 &
      while_or_2_cse_1;
  assign and_74_nl = or_5_cse & (operator_8_false_1_acc_tmp[9]);
  assign and_75_nl = or_5_cse & (~ (operator_8_false_1_acc_tmp[9]));
  assign while_while_last_burst_lpi_1_dfm_2_mx0 = MUX1HOT_s_1_3_2(while_while_if_1_if_while_while_if_1_if_nor_mx1w0,
      (~ operator_32_false_acc_itm_28_1), while_while_last_burst_lpi_1_dfm_2, {and_74_nl
      , and_75_nl , and_dcpl_14});
  assign exit_while_while_lpi_1_dfm_1_mx0w0 = while_while_last_burst_lpi_1_dfm_2_mx0
      & while_while_while_last_sva_mx1w0;
  assign while_while_while_while_or_tmp = exitL_exit_while_while_while_lpi_1 | exit_while_while_lpi_1_dfm_1
      | exitL_exit_while_while_sva;
  assign nl_operator_32_false_acc_nl = ({1'b1 , (~ while_ex_ex_len_lpi_1_dfm_31_4_mx0)})
      + 29'b00000000000000000000000000001;
  assign operator_32_false_acc_nl = nl_operator_32_false_acc_nl[28:0];
  assign operator_32_false_acc_itm_28_1 = readslicef_29_1_28(operator_32_false_acc_nl);
  assign while_while_aw_len_and_nl = (~ while_stage_v_1) & and_dcpl_14;
  assign while_while_aw_len_and_1_nl = while_stage_v_1 & and_dcpl_14;
  assign while_while_aw_len_lpi_1_dfm_3_mx0 = MUX1HOT_v_8_3_2(({{3{while_while_if_1_mux_2_psp_mx0[4]}},
      while_while_if_1_mux_2_psp_mx0}), while_while_aw_len_lpi_1, while_while_aw_len_sva_4,
      {(~ and_dcpl_14) , while_while_aw_len_and_nl , while_while_aw_len_and_1_nl});
  assign nl_while_while_aw_len_sva_2_4_0_2 = ({1'b1 , (~ (operator_8_false_1_acc_tmp[3:0]))})
      + conv_u2u_4_5(while_while_while_while_or_3_psp_1) + 5'b00001;
  assign while_while_aw_len_sva_2_4_0_2 = nl_while_while_aw_len_sva_2_4_0_2[4:0];
  assign while_while_while_while_or_3_psp_1 = MUX_v_4_2_2(while_ex_ex_len_lpi_1_dfm_3_0_mx0,
      4'b1111, operator_32_false_acc_itm_28_1);
  assign nand_25_nl = ~((~((operator_8_false_1_acc_tmp[3:0]==4'b0000))) & (operator_8_false_1_acc_tmp[9]));
  assign while_while_if_1_mux_2_psp_mx0 = MUX_v_5_2_2(while_while_aw_len_sva_2_4_0_2,
      ({1'b0 , while_while_while_while_or_3_psp_1}), nand_25_nl);
  assign nl_operator_8_false_1_acc_tmp = conv_u2u_9_10({(while_ex_addr_31_3_lpi_1_dfm_28_4_mx0[4:0])
      , while_ex_addr_31_3_lpi_1_dfm_3_0_mx0}) + conv_u2u_4_10(while_while_while_while_or_3_psp_1)
      + 10'b0000000001;
  assign operator_8_false_1_acc_tmp = nl_operator_8_false_1_acc_tmp[9:0];
  assign while_ex_addr_31_3_lpi_1_dfm_28_4_mx0 = MUX_v_25_2_2(while_ex_addr_31_3_lpi_1_28_4,
      (ex_aw_chan_Pop_mioi_idat_mxwt[35:11]), exitL_exit_while_while_sva);
  assign while_ex_addr_31_3_lpi_1_dfm_3_0_mx0 = MUX_v_4_2_2(while_ex_addr_31_3_lpi_1_3_0,
      (ex_aw_chan_Pop_mioi_idat_mxwt[10:7]), exitL_exit_while_while_sva);
  assign while_ex_ex_len_lpi_1_dfm_3_0_mx0 = MUX_v_4_2_2(while_ex_ex_len_lpi_1_3_0,
      (ex_aw_chan_Pop_mioi_idat_mxwt[39:36]), exitL_exit_while_while_sva);
  assign while_ex_ex_len_lpi_1_dfm_31_4_mx0 = MUX_v_28_2_2(while_ex_ex_len_lpi_1_31_4,
      (ex_aw_chan_Pop_mioi_idat_mxwt[67:40]), exitL_exit_while_while_sva);
  assign nl_while_while_aw_len_sva_4 = while_while_aw_len_lpi_1 + 8'b11111111;
  assign while_while_aw_len_sva_4 = nl_while_while_aw_len_sva_4[7:0];
  assign while_or_cse_1 = aw_out_Push_mioi_bawt | (~(exitL_exit_while_while_while_lpi_1_dfm_st_1
      & while_stage_v_1));
  assign while_or_1_cse_1 = last_bit_chan_Push_mioi_bawt | (~ while_stage_v_1);
  assign while_or_2_cse_1 = last_burst_chan_Push_mioi_bawt | (~(while_while_while_last_sva_st_1
      & while_stage_v_1));
  assign while_while_mux_13_nl = MUX_v_25_2_2((z_out[28:4]), (z_out[24:0]), operator_32_false_acc_itm_28_1);
  assign while_while_mux_12_nl = MUX_v_4_2_2((z_out[3:0]), while_ex_addr_31_3_lpi_1_dfm_3_0_mx0,
      operator_32_false_acc_itm_28_1);
  assign nl_while_ex_addr_31_3_sva_5 = ({while_while_mux_13_nl , while_while_mux_12_nl})
      + conv_s2u_5_29({1'b1 , (~ (operator_8_false_1_acc_tmp[3:0]))}) + 29'b00000000000000000000000000001;
  assign while_ex_addr_31_3_sva_5 = nl_while_ex_addr_31_3_sva_5[28:0];
  assign nl_while_ex_ex_len_sva_4 = ({while_ex_ex_len_lpi_1_dfm_1_31_4_1 , while_ex_ex_len_lpi_1_dfm_1_3_0_1})
      + conv_u2u_4_32(operator_8_false_1_acc_tmp[3:0]);
  assign while_ex_ex_len_sva_4 = nl_while_ex_ex_len_sva_4[31:0];
  assign nl_operator_32_false_acc_nl_1 = while_ex_ex_len_lpi_1_dfm_31_4_mx0 + 28'b1111111111111111111111111111;
  assign operator_32_false_acc_nl_1 = nl_operator_32_false_acc_nl_1[27:0];
  assign while_while_not_26_nl = ~ operator_32_false_acc_itm_28_1;
  assign while_ex_ex_len_lpi_1_dfm_1_31_4_1 = MUX_v_28_2_2(operator_32_false_acc_nl_1,
      28'b1111111111111111111111111111, while_while_not_26_nl);
  assign while_while_not_22_nl = ~ operator_32_false_acc_itm_28_1;
  assign while_ex_ex_len_lpi_1_dfm_1_3_0_1 = MUX_v_4_2_2(while_ex_ex_len_lpi_1_dfm_3_0_mx0,
      4'b1111, while_while_not_22_nl);
  assign while_while_while_asn_12 = and_137_cse & while_while_while_while_or_tmp;
  assign while_while_if_1_mux_2_tmp = MUX_v_5_2_2(({1'b0 , while_while_while_while_or_3_psp_1}),
      while_while_aw_len_sva_2_4_0_2, and_137_cse);
  assign or_dcpl_4 = exitL_exit_while_while_while_lpi_1 | exit_while_while_lpi_1_dfm_1;
  assign or_5_cse = or_dcpl_4 | exitL_exit_while_while_sva;
  assign or_19_cse = aw_out_Push_mioi_bawt | (~ exitL_exit_while_while_while_lpi_1_dfm_st_1);
  assign nand_tmp_6 = ~(while_while_last_burst_lpi_1_dfm_2 & mux_30_cse);
  assign and_dcpl_4 = while_while_asn_itm & (~ ex_aw_chan_Pop_mioi_bawt);
  assign and_dcpl_7 = or_106_cse & while_stage_v_1;
  assign or_dcpl_21 = and_dcpl_7 | and_dcpl_4;
  assign and_dcpl_14 = ~(exitL_exit_while_while_while_lpi_1 | exit_while_while_lpi_1_dfm_1
      | exitL_exit_while_while_sva);
  assign and_dcpl_15 = while_while_aw_out_write_reset_check_ResetChecker_nand_cse
      & or_49_cse;
  assign and_dcpl_18 = and_dcpl_15 & or_dcpl_4 & (~ exitL_exit_while_while_sva);
  assign and_dcpl_19 = ~((while_while_if_1_mux_2_tmp[4:3]!=2'b00));
  assign and_dcpl_22 = ~((while_while_if_1_mux_2_tmp[2:0]!=3'b000));
  assign and_dcpl_24 = and_dcpl_15 & or_5_cse;
  assign and_dcpl_37 = or_19_cse & or_132_cse;
  assign or_tmp_78 = and_dcpl_15 & (fsm_output[1]);
  assign while_stage_v_1_mx0c1 = and_dcpl_37 & last_bit_chan_Push_mioi_bawt & while_while_asn_itm
      & (~ ex_aw_chan_Pop_mioi_bawt) & while_stage_v_1;
  assign or_tmp_92 = operator_32_false_acc_itm_28_1 & (fsm_output[1]);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_aw_chan_Pop_mioi_iswt0 <= 1'b0;
      last_burst_chan_Push_mioi_m_rsc_dat <= 1'b0;
      last_burst_chan_Push_mioi_iswt0 <= 1'b0;
      last_bit_chan_Push_mioi_m_rsc_dat <= 1'b0;
      last_bit_chan_Push_mioi_iswt0 <= 1'b0;
      aw_out_Push_mioi_iswt0 <= 1'b0;
      while_while_last_burst_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( ex_aw_process_wen ) begin
      ex_aw_chan_Pop_mioi_iswt0 <= ~((mux_29_nl | (~ while_stage_en_1_mx0w1)) & (fsm_output[1]));
      last_burst_chan_Push_mioi_m_rsc_dat <= while_while_mux_5_rmff;
      last_burst_chan_Push_mioi_iswt0 <= and_103_rmff;
      last_bit_chan_Push_mioi_m_rsc_dat <= while_while_while_mux_rmff;
      last_bit_chan_Push_mioi_iswt0 <= or_tmp_78;
      aw_out_Push_mioi_iswt0 <= and_dcpl_24 & (fsm_output[1]);
      while_while_last_burst_lpi_1_dfm_2 <= while_while_last_burst_lpi_1_dfm_2_mx0;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      exitL_exit_while_while_sva <= 1'b1;
      exit_while_while_lpi_1_dfm_1 <= 1'b0;
      while_while_while_last_sva_st_1 <= 1'b0;
      exitL_exit_while_while_while_lpi_1_dfm_st_1 <= 1'b0;
    end
    else if ( while_while_and_cse ) begin
      exitL_exit_while_while_sva <= exit_while_while_lpi_1_dfm_1_mx0w0;
      exit_while_while_lpi_1_dfm_1 <= exit_while_while_lpi_1_dfm_1_mx0w0;
      while_while_while_last_sva_st_1 <= while_while_while_last_sva_mx1w0;
      exitL_exit_while_while_while_lpi_1_dfm_st_1 <= while_while_while_while_or_tmp;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      aw_out_Push_mioi_idat_40_36 <= 5'b00000;
    end
    else if ( while_while_and_1_cse & ((or_56_cse & while_while_aw_out_write_reset_check_ResetChecker_nand_cse
        & or_49_cse & or_5_cse & (operator_8_false_1_acc_tmp[9])) | and_28_rgt) )
        begin
      aw_out_Push_mioi_idat_40_36 <= MUX_v_5_2_2(while_while_aw_len_sva_2_4_0_2,
          ({1'b0 , while_while_while_while_or_3_psp_1}), and_28_rgt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      aw_out_Push_mioi_idat_10_7 <= 4'b0000;
      aw_out_Push_mioi_idat_35_11 <= 25'b0000000000000000000000000;
      aw_out_Push_mioi_idat_6_0 <= 7'b0000000;
    end
    else if ( while_while_and_9_cse ) begin
      aw_out_Push_mioi_idat_10_7 <= MUX_v_4_2_2((ex_aw_chan_Pop_mioi_idat_mxwt[10:7]),
          while_ex_addr_31_3_lpi_1_3_0, and_dcpl_18);
      aw_out_Push_mioi_idat_35_11 <= MUX_v_25_2_2((ex_aw_chan_Pop_mioi_idat_mxwt[35:11]),
          while_ex_addr_31_3_lpi_1_28_4, and_dcpl_18);
      aw_out_Push_mioi_idat_6_0 <= MUX_v_7_2_2((ex_aw_chan_Pop_mioi_idat_mxwt[6:0]),
          assocmrg_lpi_1_dfm_6_0, and_dcpl_18);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_while_asn_itm <= 1'b1;
    end
    else if ( ex_aw_process_wen & ((while_stage_en_1_mx0w1 & (fsm_output[1])) | ((~
        while_while_asn_itm) & while_stage_en_1_mx0w1)) ) begin
      while_while_asn_itm <= exit_while_while_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      assocmrg_lpi_1_dfm_6_0 <= 7'b0000000;
    end
    else if ( ex_aw_process_wen & exitL_exit_while_while_sva ) begin
      assocmrg_lpi_1_dfm_6_0 <= ex_aw_chan_Pop_mioi_idat_mxwt[6:0];
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_while_aw_len_lpi_1 <= 8'b00000000;
    end
    else if ( ex_aw_process_wen & ((and_15_cse & and_dcpl_4 & while_stage_v_1) |
        (while_stage_v_1 & and_15_cse & or_49_cse & and_dcpl_14) | and_78_rgt) )
        begin
      while_while_aw_len_lpi_1 <= MUX_v_8_2_2(while_while_aw_len_sva_4, ({{3{while_while_if_1_mux_2_psp_mx0[4]}},
          while_while_if_1_mux_2_psp_mx0}), and_78_rgt);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_ex_addr_31_3_lpi_1_28_4 <= 25'b0000000000000000000000000;
      while_ex_ex_len_lpi_1_31_4 <= 28'b0000000000000000000000000000;
      while_ex_ex_len_lpi_1_3_0 <= 4'b0000;
    end
    else if ( while_ex_addr_and_cse ) begin
      while_ex_addr_31_3_lpi_1_28_4 <= MUX_v_25_2_2((z_out[24:0]), (while_ex_addr_31_3_sva_5[28:4]),
          while_ex_addr_and_4_cse);
      while_ex_ex_len_lpi_1_31_4 <= MUX_v_28_2_2(while_ex_ex_len_lpi_1_dfm_1_31_4_1,
          (while_ex_ex_len_sva_4[31:4]), while_ex_addr_and_4_cse);
      while_ex_ex_len_lpi_1_3_0 <= MUX_v_4_2_2(while_ex_ex_len_lpi_1_dfm_1_3_0_1,
          (while_ex_ex_len_sva_4[3:0]), while_ex_addr_and_4_cse);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_ex_addr_31_3_lpi_1_3_0 <= 4'b0000;
    end
    else if ( ex_aw_process_wen & ((exitL_exit_while_while_sva & (~(while_while_while_asn_12
        | or_dcpl_21))) | while_ex_addr_and_4_cse) ) begin
      while_ex_addr_31_3_lpi_1_3_0 <= MUX_v_4_2_2((ex_aw_chan_Pop_mioi_idat_mxwt[10:7]),
          (while_ex_addr_31_3_sva_5[3:0]), while_ex_addr_and_4_cse);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      exitL_exit_while_while_while_lpi_1 <= 1'b0;
    end
    else if ( ex_aw_process_wen & (~ or_dcpl_21) ) begin
      exitL_exit_while_while_while_lpi_1 <= while_while_while_last_sva_mx1w0;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_stage_v_1 <= 1'b0;
    end
    else if ( ex_aw_process_wen & (or_tmp_78 | while_stage_v_1_mx0c1) ) begin
      while_stage_v_1 <= ~ while_stage_v_1_mx0c1;
    end
  end
  assign mux_26_nl = MUX_s_1_2_2((~ nand_tmp_6), nand_1_cse, or_dcpl_4);
  assign nor_10_nl = ~(exitL_exit_while_while_sva | mux_26_nl);
  assign or_58_nl = (operator_8_false_1_acc_tmp[9]) | (~ nand_1_cse);
  assign mux_24_nl = MUX_s_1_2_2(nand_tmp_6, or_58_nl, or_dcpl_4);
  assign and_18_nl = (operator_8_false_1_acc_tmp[9]) & nand_1_cse;
  assign mux_25_nl = MUX_s_1_2_2(mux_24_nl, and_18_nl, exitL_exit_while_while_sva);
  assign mux_27_nl = MUX_s_1_2_2(nor_10_nl, mux_25_nl, or_56_cse);
  assign nand_5_nl = ~((~(exit_while_while_lpi_1_dfm_1 | exitL_exit_while_while_while_lpi_1
      | (~ while_while_last_burst_lpi_1_dfm_2))) & mux_30_cse);
  assign mux_23_nl = MUX_s_1_2_2(nand_5_nl, nand_1_cse, exitL_exit_while_while_sva);
  assign or_50_nl = (while_while_if_1_mux_2_tmp!=5'b00000) | operator_32_false_acc_itm_28_1;
  assign mux_28_nl = MUX_s_1_2_2(mux_27_nl, mux_23_nl, or_50_nl);
  assign mux_29_nl = MUX_s_1_2_2((~ exitL_exit_while_while_sva), mux_28_nl, or_49_cse);
  assign operator_8_false_mux_2_nl = MUX_v_29_2_2(({while_ex_addr_31_3_lpi_1_dfm_28_4_mx0
      , while_ex_addr_31_3_lpi_1_dfm_3_0_mx0}), ({4'b0000 , while_ex_addr_31_3_lpi_1_dfm_28_4_mx0}),
      or_tmp_92);
  assign operator_8_false_operator_8_false_nand_1_nl = ~(or_tmp_92 & (~((~ operator_32_false_acc_itm_28_1)
      & (fsm_output[1]))));
  assign operator_8_false_mux_3_nl = MUX_v_4_2_2(while_ex_ex_len_lpi_1_dfm_3_0_mx0,
      4'b0001, or_tmp_92);
  assign nl_acc_nl = ({operator_8_false_mux_2_nl , operator_8_false_operator_8_false_nand_1_nl})
      + conv_u2u_5_30({operator_8_false_mux_3_nl , 1'b1});
  assign acc_nl = nl_acc_nl[29:0];
  assign z_out = readslicef_30_29_1(acc_nl);

  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & {1{sel}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & {1{sel}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input  sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [27:0] MUX_v_28_2_2;
    input [27:0] input_0;
    input [27:0] input_1;
    input  sel;
    reg [27:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_28_2_2 = result;
  end
  endfunction


  function automatic [28:0] MUX_v_29_2_2;
    input [28:0] input_0;
    input [28:0] input_1;
    input  sel;
    reg [28:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_29_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_29_1_28;
    input [28:0] vector;
    reg [28:0] tmp;
  begin
    tmp = vector >> 28;
    readslicef_29_1_28 = tmp[0:0];
  end
  endfunction


  function automatic [28:0] readslicef_30_29_1;
    input [29:0] vector;
    reg [29:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_30_29_1 = tmp[28:0];
  end
  endfunction


  function automatic [43:0] signext_44_41;
    input [40:0] vector;
  begin
    signext_44_41= {{3{vector[40]}}, vector};
  end
  endfunction


  function automatic [28:0] conv_s2u_5_29 ;
    input [4:0]  vector ;
  begin
    conv_s2u_5_29 = {{24{vector[4]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_4_10 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_10 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_4_32 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_32 = {{28{1'b0}}, vector};
  end
  endfunction


  function automatic [29:0] conv_u2u_5_30 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_30 = {{25{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process (
  clk, rst_bar, ar_out_vld, ar_out_rdy, ar_out_dat, ex_ar_chan_vld, ex_ar_chan_rdy,
      ex_ar_chan_dat
);
  input clk;
  input rst_bar;
  output ar_out_vld;
  input ar_out_rdy;
  output [43:0] ar_out_dat;
  input ex_ar_chan_vld;
  output ex_ar_chan_rdy;
  input [75:0] ex_ar_chan_dat;


  // Interconnect Declarations
  wire ex_ar_process_wen;
  wire ex_ar_process_wten;
  wire ex_ar_chan_Pop_mioi_bawt;
  reg ex_ar_chan_Pop_mioi_iswt0;
  wire ex_ar_chan_Pop_mioi_wen_comp;
  wire [67:0] ex_ar_chan_Pop_mioi_idat_mxwt;
  wire ar_out_Push_mioi_bawt;
  reg ar_out_Push_mioi_iswt0;
  wire ar_out_Push_mioi_wen_comp;
  reg [6:0] ar_out_Push_mioi_idat_6_0;
  reg [24:0] ar_out_Push_mioi_idat_35_11;
  reg [3:0] ar_out_Push_mioi_idat_10_7;
  reg [4:0] ar_out_Push_mioi_idat_40_36;
  wire [1:0] fsm_output;
  wire [9:0] operator_8_false_1_acc_tmp;
  wire [10:0] nl_operator_8_false_1_acc_tmp;
  wire nand_tmp;
  wire and_dcpl_3;
  wire and_dcpl_10;
  wire and_dcpl_12;
  wire and_dcpl_17;
  wire and_dcpl_18;
  wire and_dcpl_21;
  wire and_dcpl_22;
  wire and_dcpl_25;
  wire and_dcpl_27;
  wire and_dcpl_29;
  wire or_dcpl_14;
  wire and_dcpl_37;
  wire and_dcpl_38;
  wire and_dcpl_39;
  wire or_tmp_38;
  wire while_stage_en_1_mx0w1;
  reg while_while_asn_itm;
  reg while_stage_v_1;
  reg exitL_exit_while_while_sva;
  reg while_while_if_1_and_2_itm_1;
  wire or_66_cse;
  wire or_14_cse;
  wire or_13_cse;
  wire and_86_cse;
  wire [28:0] while_ex_addr_31_3_sva_4;
  wire [29:0] nl_while_ex_addr_31_3_sva_4;
  wire or_tmp_49;
  wire [28:0] z_out;
  reg [3:0] operator_13_false_1_operator_13_false_1_slc_while_while_if_1_endbits_10_0_1_itm_1;
  reg [24:0] while_ex_addr_31_3_lpi_1_28_4;
  reg [3:0] while_ex_addr_31_3_lpi_1_3_0;
  reg [27:0] while_ex_ex_len_lpi_1_31_4;
  reg [3:0] while_ex_ex_len_lpi_1_3_0;
  reg [6:0] assocmrg_lpi_1_dfm_6_0;
  wire while_while_if_1_if_while_while_if_1_if_nor_mx0w0;
  wire exitL_exit_while_while_sva_mx0c1;
  wire ar_out_Push_mioi_idat_40_36_mx0c1;
  wire [3:0] while_while_asn_13_mx1w1;
  wire [24:0] while_while_asn_11_mx1w1;
  wire while_while_asn_itm_mx0c1;
  wire while_stage_v_1_mx0c1;
  wire [3:0] while_while_while_while_or_2_psp_1;
  wire [24:0] while_ex_addr_31_3_lpi_1_dfm_28_4_mx0;
  wire [3:0] while_ex_addr_31_3_lpi_1_dfm_3_0_mx0;
  wire [3:0] while_ex_ex_len_lpi_1_dfm_3_0_mx0;
  wire [27:0] while_ex_ex_len_lpi_1_dfm_31_4_mx0;
  wire [31:0] while_ex_ex_len_sva_4;
  wire [32:0] nl_while_ex_ex_len_sva_4;
  wire [27:0] while_ex_ex_len_lpi_1_dfm_1_31_4_1;
  wire [3:0] while_ex_ex_len_lpi_1_dfm_1_3_0_1;
  wire while_while_and_7_cse;
  wire while_ex_addr_and_cse;
  wire while_ex_ex_len_and_cse;
  wire operator_13_false_1_and_cse;
  wire operator_32_false_acc_itm_28_1;

  wire mux_17_nl;
  wire and_nl;
  wire[4:0] while_while_if_1_if_if_acc_nl;
  wire[5:0] nl_while_while_if_1_if_if_acc_nl;
  wire[28:0] operator_32_false_acc_nl;
  wire[29:0] nl_operator_32_false_acc_nl;
  wire[27:0] operator_32_false_acc_nl_1;
  wire[28:0] nl_operator_32_false_acc_nl_1;
  wire while_while_not_20_nl;
  wire while_while_not_21_nl;
  wire[29:0] acc_nl;
  wire[30:0] nl_acc_nl;
  wire[28:0] operator_32_false_mux_2_nl;
  wire operator_32_false_or_1_nl;
  wire[3:0] operator_32_false_mux_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_inst_ex_ar_chan_Pop_mioi_oswt_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_inst_ex_ar_chan_Pop_mioi_oswt_unreg
      = or_13_cse & while_while_asn_itm & ex_ar_chan_Pop_mioi_bawt & (fsm_output[1]);
  wire [43:0] nl_axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_inst_ar_out_Push_mioi_idat;
  assign nl_axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_inst_ar_out_Push_mioi_idat
      = signext_44_41({ar_out_Push_mioi_idat_40_36 , ar_out_Push_mioi_idat_35_11
      , ar_out_Push_mioi_idat_10_7 , ar_out_Push_mioi_idat_6_0});
  wire  nl_axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_staller_inst_ex_ar_process_flen_unreg;
  assign nl_axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_staller_inst_ex_ar_process_flen_unreg
      = ~((~((~ while_stage_en_1_mx0w1) & (fsm_output[1]))) | (while_stage_en_1_mx0w1
      & (fsm_output[1])) | (while_stage_v_1 & or_13_cse & (fsm_output[1])));
  axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_ar_chan_vld(ex_ar_chan_vld),
      .ex_ar_chan_rdy(ex_ar_chan_rdy),
      .ex_ar_chan_dat(ex_ar_chan_dat),
      .ex_ar_process_wen(ex_ar_process_wen),
      .ex_ar_process_wten(ex_ar_process_wten),
      .ex_ar_chan_Pop_mioi_oswt_unreg(nl_axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_chan_Pop_mioi_inst_ex_ar_chan_Pop_mioi_oswt_unreg),
      .ex_ar_chan_Pop_mioi_bawt(ex_ar_chan_Pop_mioi_bawt),
      .ex_ar_chan_Pop_mioi_iswt0(ex_ar_chan_Pop_mioi_iswt0),
      .ex_ar_chan_Pop_mioi_wen_comp(ex_ar_chan_Pop_mioi_wen_comp),
      .ex_ar_chan_Pop_mioi_idat_mxwt(ex_ar_chan_Pop_mioi_idat_mxwt)
    );
  axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ar_out_vld(ar_out_vld),
      .ar_out_rdy(ar_out_rdy),
      .ar_out_dat(ar_out_dat),
      .ex_ar_process_wen(ex_ar_process_wen),
      .ex_ar_process_wten(ex_ar_process_wten),
      .ar_out_Push_mioi_oswt_unreg(and_dcpl_22),
      .ar_out_Push_mioi_bawt(ar_out_Push_mioi_bawt),
      .ar_out_Push_mioi_iswt0(ar_out_Push_mioi_iswt0),
      .ar_out_Push_mioi_wen_comp(ar_out_Push_mioi_wen_comp),
      .ar_out_Push_mioi_idat(nl_axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ar_out_Push_mioi_inst_ar_out_Push_mioi_idat[43:0])
    );
  axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_staller axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_staller_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_ar_process_wen(ex_ar_process_wen),
      .ex_ar_process_wten(ex_ar_process_wten),
      .ex_ar_chan_Pop_mioi_wen_comp(ex_ar_chan_Pop_mioi_wen_comp),
      .ar_out_Push_mioi_wen_comp(ar_out_Push_mioi_wen_comp),
      .ex_ar_process_flen_unreg(nl_axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_staller_inst_ex_ar_process_flen_unreg)
    );
  axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_process_fsm axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_ex_ar_process_fsm_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ex_ar_process_wen(ex_ar_process_wen),
      .fsm_output(fsm_output)
    );
  assign or_66_cse = (operator_8_false_1_acc_tmp[3:0]!=4'b0000);
  assign and_86_cse = or_66_cse & (operator_8_false_1_acc_tmp[9]);
  assign while_while_and_7_cse = ex_ar_process_wen & (~ (fsm_output[0])) & ((while_stage_en_1_mx0w1
      & exitL_exit_while_while_sva) | and_dcpl_21);
  assign while_ex_addr_and_cse = ex_ar_process_wen & (and_dcpl_37 | and_dcpl_38 |
      and_dcpl_39);
  assign while_ex_ex_len_and_cse = ex_ar_process_wen & (and_dcpl_12 | and_dcpl_18);
  assign or_14_cse = (~ while_while_asn_itm) | ex_ar_chan_Pop_mioi_bawt;
  assign or_13_cse = (~ while_stage_v_1) | ar_out_Push_mioi_bawt;
  assign operator_13_false_1_and_cse = ex_ar_process_wen & (~(while_stage_v_1 & (~
      ar_out_Push_mioi_bawt)));
  assign while_while_if_1_if_while_while_if_1_if_nor_mx0w0 = ~(operator_32_false_acc_itm_28_1
      | or_66_cse);
  assign while_while_asn_13_mx1w1 = MUX_v_4_2_2((while_ex_addr_31_3_sva_4[3:0]),
      while_ex_addr_31_3_lpi_1_3_0, or_dcpl_14);
  assign while_while_asn_11_mx1w1 = MUX_v_25_2_2((while_ex_addr_31_3_sva_4[28:4]),
      while_ex_addr_31_3_lpi_1_28_4, or_dcpl_14);
  assign while_stage_en_1_mx0w1 = or_14_cse & or_13_cse;
  assign while_while_while_while_or_2_psp_1 = MUX_v_4_2_2(while_ex_ex_len_lpi_1_dfm_3_0_mx0,
      4'b1111, operator_32_false_acc_itm_28_1);
  assign nl_operator_8_false_1_acc_tmp = conv_u2u_9_10({(while_ex_addr_31_3_lpi_1_dfm_28_4_mx0[4:0])
      , while_ex_addr_31_3_lpi_1_dfm_3_0_mx0}) + conv_u2u_4_10(while_while_while_while_or_2_psp_1)
      + 10'b0000000001;
  assign operator_8_false_1_acc_tmp = nl_operator_8_false_1_acc_tmp[9:0];
  assign nl_operator_32_false_acc_nl = ({1'b1 , (~ while_ex_ex_len_lpi_1_dfm_31_4_mx0)})
      + 29'b00000000000000000000000000001;
  assign operator_32_false_acc_nl = nl_operator_32_false_acc_nl[28:0];
  assign operator_32_false_acc_itm_28_1 = readslicef_29_1_28(operator_32_false_acc_nl);
  assign while_ex_addr_31_3_lpi_1_dfm_28_4_mx0 = MUX_v_25_2_2(while_while_asn_11_mx1w1,
      (ex_ar_chan_Pop_mioi_idat_mxwt[35:11]), exitL_exit_while_while_sva);
  assign while_ex_addr_31_3_lpi_1_dfm_3_0_mx0 = MUX_v_4_2_2(while_while_asn_13_mx1w1,
      (ex_ar_chan_Pop_mioi_idat_mxwt[10:7]), exitL_exit_while_while_sva);
  assign while_ex_ex_len_lpi_1_dfm_3_0_mx0 = MUX_v_4_2_2(while_ex_ex_len_lpi_1_3_0,
      (ex_ar_chan_Pop_mioi_idat_mxwt[39:36]), exitL_exit_while_while_sva);
  assign while_ex_ex_len_lpi_1_dfm_31_4_mx0 = MUX_v_28_2_2(while_ex_ex_len_lpi_1_31_4,
      (ex_ar_chan_Pop_mioi_idat_mxwt[67:40]), exitL_exit_while_while_sva);
  assign nl_while_ex_addr_31_3_sva_4 = ({while_ex_addr_31_3_lpi_1_28_4 , while_ex_addr_31_3_lpi_1_3_0})
      + conv_s2u_5_29({1'b1 , (~ operator_13_false_1_operator_13_false_1_slc_while_while_if_1_endbits_10_0_1_itm_1)})
      + 29'b00000000000000000000000000001;
  assign while_ex_addr_31_3_sva_4 = nl_while_ex_addr_31_3_sva_4[28:0];
  assign nl_while_ex_ex_len_sva_4 = ({while_ex_ex_len_lpi_1_dfm_1_31_4_1 , while_ex_ex_len_lpi_1_dfm_1_3_0_1})
      + conv_u2u_4_32(operator_8_false_1_acc_tmp[3:0]);
  assign while_ex_ex_len_sva_4 = nl_while_ex_ex_len_sva_4[31:0];
  assign nl_operator_32_false_acc_nl_1 = while_ex_ex_len_lpi_1_dfm_31_4_mx0 + 28'b1111111111111111111111111111;
  assign operator_32_false_acc_nl_1 = nl_operator_32_false_acc_nl_1[27:0];
  assign while_while_not_20_nl = ~ operator_32_false_acc_itm_28_1;
  assign while_ex_ex_len_lpi_1_dfm_1_31_4_1 = MUX_v_28_2_2(operator_32_false_acc_nl_1,
      28'b1111111111111111111111111111, while_while_not_20_nl);
  assign while_while_not_21_nl = ~ operator_32_false_acc_itm_28_1;
  assign while_ex_ex_len_lpi_1_dfm_1_3_0_1 = MUX_v_4_2_2(while_ex_ex_len_lpi_1_dfm_3_0_mx0,
      4'b1111, while_while_not_21_nl);
  assign nand_tmp = ~(exitL_exit_while_while_sva & (~ while_stage_en_1_mx0w1));
  assign and_dcpl_3 = (~ while_while_asn_itm) & (operator_8_false_1_acc_tmp[9]);
  assign and_dcpl_10 = or_66_cse & or_13_cse;
  assign and_dcpl_12 = and_dcpl_10 & or_14_cse & (operator_8_false_1_acc_tmp[9]);
  assign and_dcpl_17 = (~((~((operator_8_false_1_acc_tmp[3:0]==4'b0000))) & (operator_8_false_1_acc_tmp[9])))
      & or_13_cse;
  assign and_dcpl_18 = and_dcpl_17 & or_14_cse;
  assign and_dcpl_21 = while_stage_en_1_mx0w1 & (~ exitL_exit_while_while_sva);
  assign and_dcpl_22 = while_stage_v_1 & ar_out_Push_mioi_bawt;
  assign and_dcpl_25 = (operator_8_false_1_acc_tmp[9]) & while_stage_en_1_mx0w1;
  assign and_dcpl_27 = or_13_cse & (~ while_while_asn_itm);
  assign and_dcpl_29 = (~ (operator_8_false_1_acc_tmp[9])) & while_stage_en_1_mx0w1;
  assign or_dcpl_14 = ~(while_stage_v_1 & while_while_if_1_and_2_itm_1);
  assign and_dcpl_37 = and_dcpl_22 & while_while_asn_itm & (~ ex_ar_chan_Pop_mioi_bawt)
      & while_while_if_1_and_2_itm_1;
  assign and_dcpl_38 = while_stage_en_1_mx0w1 & operator_32_false_acc_itm_28_1;
  assign and_dcpl_39 = while_stage_en_1_mx0w1 & (~ operator_32_false_acc_itm_28_1);
  assign or_tmp_38 = while_stage_en_1_mx0w1 & (fsm_output[1]);
  assign exitL_exit_while_while_sva_mx0c1 = (while_stage_en_1_mx0w1 & (~ (operator_8_false_1_acc_tmp[9]))
      & (fsm_output[1])) | (or_13_cse & (~ while_while_asn_itm) & (~ (operator_8_false_1_acc_tmp[9])));
  assign ar_out_Push_mioi_idat_40_36_mx0c1 = (and_dcpl_18 & (fsm_output[1])) | (and_dcpl_17
      & (~ while_while_asn_itm));
  assign while_while_asn_itm_mx0c1 = (and_dcpl_29 & (fsm_output[1])) | (and_dcpl_27
      & and_dcpl_29);
  assign while_stage_v_1_mx0c1 = and_dcpl_22 & while_while_asn_itm & (~ ex_ar_chan_Pop_mioi_bawt);
  assign or_tmp_49 = (~ operator_32_false_acc_itm_28_1) & (fsm_output[1]);
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ex_ar_chan_Pop_mioi_iswt0 <= 1'b0;
      ar_out_Push_mioi_iswt0 <= 1'b0;
    end
    else if ( ex_ar_process_wen ) begin
      ex_ar_chan_Pop_mioi_iswt0 <= ~((mux_17_nl | (~ while_stage_en_1_mx0w1)) & (fsm_output[1]));
      ar_out_Push_mioi_iswt0 <= or_tmp_38;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      exitL_exit_while_while_sva <= 1'b1;
    end
    else if ( ex_ar_process_wen & ((while_stage_en_1_mx0w1 & (operator_8_false_1_acc_tmp[9])
        & (fsm_output[1])) | (or_13_cse & and_dcpl_3) | exitL_exit_while_while_sva_mx0c1)
        ) begin
      exitL_exit_while_while_sva <= MUX_s_1_2_2(while_while_if_1_if_while_while_if_1_if_nor_mx0w0,
          (~ operator_32_false_acc_itm_28_1), exitL_exit_while_while_sva_mx0c1);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ar_out_Push_mioi_idat_40_36 <= 5'b00000;
    end
    else if ( ex_ar_process_wen & ((and_dcpl_12 & (fsm_output[1])) | (and_dcpl_10
        & and_dcpl_3) | ar_out_Push_mioi_idat_40_36_mx0c1) ) begin
      ar_out_Push_mioi_idat_40_36 <= MUX_v_5_2_2(while_while_if_1_if_if_acc_nl, ({1'b0
          , while_while_while_while_or_2_psp_1}), ar_out_Push_mioi_idat_40_36_mx0c1);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      ar_out_Push_mioi_idat_10_7 <= 4'b0000;
      ar_out_Push_mioi_idat_35_11 <= 25'b0000000000000000000000000;
      ar_out_Push_mioi_idat_6_0 <= 7'b0000000;
    end
    else if ( while_while_and_7_cse ) begin
      ar_out_Push_mioi_idat_10_7 <= MUX_v_4_2_2((ex_ar_chan_Pop_mioi_idat_mxwt[10:7]),
          while_while_asn_13_mx1w1, and_dcpl_21);
      ar_out_Push_mioi_idat_35_11 <= MUX_v_25_2_2((ex_ar_chan_Pop_mioi_idat_mxwt[35:11]),
          while_while_asn_11_mx1w1, and_dcpl_21);
      ar_out_Push_mioi_idat_6_0 <= MUX_v_7_2_2((ex_ar_chan_Pop_mioi_idat_mxwt[6:0]),
          assocmrg_lpi_1_dfm_6_0, and_dcpl_21);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_while_asn_itm <= 1'b1;
    end
    else if ( ex_ar_process_wen & ((and_dcpl_25 & (fsm_output[1])) | (and_dcpl_27
        & and_dcpl_25) | while_while_asn_itm_mx0c1) ) begin
      while_while_asn_itm <= MUX_s_1_2_2(while_while_if_1_if_while_while_if_1_if_nor_mx0w0,
          (~ operator_32_false_acc_itm_28_1), while_while_asn_itm_mx0c1);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_ex_addr_31_3_lpi_1_28_4 <= 25'b0000000000000000000000000;
      while_ex_addr_31_3_lpi_1_3_0 <= 4'b0000;
    end
    else if ( while_ex_addr_and_cse ) begin
      while_ex_addr_31_3_lpi_1_28_4 <= MUX1HOT_v_25_3_2((while_ex_addr_31_3_sva_4[28:4]),
          (z_out[24:0]), (z_out[28:4]), {and_dcpl_37 , and_dcpl_38 , and_dcpl_39});
      while_ex_addr_31_3_lpi_1_3_0 <= MUX1HOT_v_4_3_2((while_ex_addr_31_3_sva_4[3:0]),
          while_ex_addr_31_3_lpi_1_dfm_3_0_mx0, (z_out[3:0]), {and_dcpl_37 , and_dcpl_38
          , and_dcpl_39});
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_ex_ex_len_lpi_1_31_4 <= 28'b0000000000000000000000000000;
      while_ex_ex_len_lpi_1_3_0 <= 4'b0000;
    end
    else if ( while_ex_ex_len_and_cse ) begin
      while_ex_ex_len_lpi_1_31_4 <= MUX_v_28_2_2((while_ex_ex_len_sva_4[31:4]), while_ex_ex_len_lpi_1_dfm_1_31_4_1,
          and_dcpl_18);
      while_ex_ex_len_lpi_1_3_0 <= MUX_v_4_2_2((while_ex_ex_len_sva_4[3:0]), while_ex_ex_len_lpi_1_dfm_1_3_0_1,
          and_dcpl_18);
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      assocmrg_lpi_1_dfm_6_0 <= 7'b0000000;
    end
    else if ( ex_ar_process_wen & exitL_exit_while_while_sva ) begin
      assocmrg_lpi_1_dfm_6_0 <= ex_ar_chan_Pop_mioi_idat_mxwt[6:0];
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      while_stage_v_1 <= 1'b0;
    end
    else if ( ex_ar_process_wen & (or_tmp_38 | while_stage_v_1_mx0c1) ) begin
      while_stage_v_1 <= ~ while_stage_v_1_mx0c1;
    end
  end
  always @(posedge clk or negedge rst_bar) begin
    if ( ~ rst_bar ) begin
      operator_13_false_1_operator_13_false_1_slc_while_while_if_1_endbits_10_0_1_itm_1
          <= 4'b0000;
      while_while_if_1_and_2_itm_1 <= 1'b0;
    end
    else if ( operator_13_false_1_and_cse ) begin
      operator_13_false_1_operator_13_false_1_slc_while_while_if_1_endbits_10_0_1_itm_1
          <= operator_8_false_1_acc_tmp[3:0];
      while_while_if_1_and_2_itm_1 <= and_86_cse;
    end
  end
  assign and_nl = nand_tmp & and_86_cse;
  assign mux_17_nl = MUX_s_1_2_2(and_nl, nand_tmp, operator_32_false_acc_itm_28_1);
  assign nl_while_while_if_1_if_if_acc_nl = ({1'b1 , (~ (operator_8_false_1_acc_tmp[3:0]))})
      + conv_u2s_4_5(while_while_while_while_or_2_psp_1) + 5'b00001;
  assign while_while_if_1_if_if_acc_nl = nl_while_while_if_1_if_if_acc_nl[4:0];
  assign operator_32_false_mux_2_nl = MUX_v_29_2_2(({4'b0000 , while_ex_addr_31_3_lpi_1_dfm_28_4_mx0}),
      ({while_ex_addr_31_3_lpi_1_dfm_28_4_mx0 , while_ex_addr_31_3_lpi_1_dfm_3_0_mx0}),
      or_tmp_49);
  assign operator_32_false_or_1_nl = (~(operator_32_false_acc_itm_28_1 & (fsm_output[1])))
      | or_tmp_49;
  assign operator_32_false_mux_3_nl = MUX_v_4_2_2(4'b0001, while_ex_ex_len_lpi_1_dfm_3_0_mx0,
      or_tmp_49);
  assign nl_acc_nl = ({operator_32_false_mux_2_nl , operator_32_false_or_1_nl}) +
      conv_u2u_5_30({operator_32_false_mux_3_nl , 1'b1});
  assign acc_nl = nl_acc_nl[29:0];
  assign z_out = readslicef_30_29_1(acc_nl);

  function automatic [24:0] MUX1HOT_v_25_3_2;
    input [24:0] input_2;
    input [24:0] input_1;
    input [24:0] input_0;
    input [2:0] sel;
    reg [24:0] result;
  begin
    result = input_0 & {25{sel[0]}};
    result = result | ( input_1 & {25{sel[1]}});
    result = result | ( input_2 & {25{sel[2]}});
    MUX1HOT_v_25_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input  sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [27:0] MUX_v_28_2_2;
    input [27:0] input_0;
    input [27:0] input_1;
    input  sel;
    reg [27:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_28_2_2 = result;
  end
  endfunction


  function automatic [28:0] MUX_v_29_2_2;
    input [28:0] input_0;
    input [28:0] input_1;
    input  sel;
    reg [28:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_29_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_29_1_28;
    input [28:0] vector;
    reg [28:0] tmp;
  begin
    tmp = vector >> 28;
    readslicef_29_1_28 = tmp[0:0];
  end
  endfunction


  function automatic [28:0] readslicef_30_29_1;
    input [29:0] vector;
    reg [29:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_30_29_1 = tmp[28:0];
  end
  endfunction


  function automatic [43:0] signext_44_41;
    input [40:0] vector;
  begin
    signext_44_41= {{3{vector[40]}}, vector};
  end
  endfunction


  function automatic [28:0] conv_s2u_5_29 ;
    input [4:0]  vector ;
  begin
    conv_s2u_5_29 = {{24{vector[4]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_4_10 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_10 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_4_32 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_32 = {{28{1'b0}}, vector};
  end
  endfunction


  function automatic [29:0] conv_u2u_5_30 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_30 = {{25{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_w_segment
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_w_segment (
  clk, rst_bar, aw_out_vld, aw_out_rdy, aw_out_dat, w_out_vld, w_out_rdy, w_out_dat,
      b_in_vld, b_in_rdy, b_in_dat, ex_aw_chan_vld, ex_aw_chan_rdy, ex_aw_chan_dat,
      w_chan_vld, w_chan_rdy, w_chan_dat, b_chan_vld, b_chan_rdy, b_chan_dat
);
  input clk;
  input rst_bar;
  output aw_out_vld;
  input aw_out_rdy;
  output [43:0] aw_out_dat;
  output w_out_vld;
  input w_out_rdy;
  output [72:0] w_out_dat;
  input b_in_vld;
  output b_in_rdy;
  input [5:0] b_in_dat;
  input ex_aw_chan_vld;
  output ex_aw_chan_rdy;
  input [75:0] ex_aw_chan_dat;
  input w_chan_vld;
  output w_chan_rdy;
  input [72:0] w_chan_dat;
  output b_chan_vld;
  input b_chan_rdy;
  output [5:0] b_chan_dat;


  // Interconnect Declarations
  wire last_bit_chan_vld;
  wire last_bit_chan_rdy;
  wire last_bit_chan_dat;
  wire last_burst_chan_vld;
  wire last_burst_chan_rdy;
  wire last_burst_chan_dat;


  // Interconnect Declarations for Component Instantiations 
  axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process axi_axi4_segment_axi_cfg_standard_w_segment_ex_aw_process_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .aw_out_vld(aw_out_vld),
      .aw_out_rdy(aw_out_rdy),
      .aw_out_dat(aw_out_dat),
      .ex_aw_chan_vld(ex_aw_chan_vld),
      .ex_aw_chan_rdy(ex_aw_chan_rdy),
      .ex_aw_chan_dat(ex_aw_chan_dat),
      .last_bit_chan_vld(last_bit_chan_vld),
      .last_bit_chan_rdy(last_bit_chan_rdy),
      .last_bit_chan_dat(last_bit_chan_dat),
      .last_burst_chan_vld(last_burst_chan_vld),
      .last_burst_chan_rdy(last_burst_chan_rdy),
      .last_burst_chan_dat(last_burst_chan_dat)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_w_process axi_axi4_segment_axi_cfg_standard_w_segment_w_process_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_out_vld(w_out_vld),
      .w_out_rdy(w_out_rdy),
      .w_out_dat(w_out_dat),
      .w_chan_vld(w_chan_vld),
      .w_chan_rdy(w_chan_rdy),
      .w_chan_dat(w_chan_dat),
      .last_bit_chan_vld(last_bit_chan_vld),
      .last_bit_chan_rdy(last_bit_chan_rdy),
      .last_bit_chan_dat(last_bit_chan_dat)
    );
  axi_axi4_segment_axi_cfg_standard_w_segment_b_process axi_axi4_segment_axi_cfg_standard_w_segment_b_process_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .b_in_vld(b_in_vld),
      .b_in_rdy(b_in_rdy),
      .b_in_dat(b_in_dat),
      .b_chan_vld(b_chan_vld),
      .b_chan_rdy(b_chan_rdy),
      .b_chan_dat(b_chan_dat),
      .last_burst_chan_vld(last_burst_chan_vld),
      .last_burst_chan_rdy(last_burst_chan_rdy),
      .last_burst_chan_dat(last_burst_chan_dat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    axi_axi4_segment_axi_cfg_standard_r_segment
// ------------------------------------------------------------------


module axi_axi4_segment_axi_cfg_standard_r_segment (
  clk, rst_bar, ar_out_vld, ar_out_rdy, ar_out_dat, ex_ar_chan_vld, ex_ar_chan_rdy,
      ex_ar_chan_dat
);
  input clk;
  input rst_bar;
  output ar_out_vld;
  input ar_out_rdy;
  output [43:0] ar_out_dat;
  input ex_ar_chan_vld;
  output ex_ar_chan_rdy;
  input [75:0] ex_ar_chan_dat;



  // Interconnect Declarations for Component Instantiations 
  axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process axi_axi4_segment_axi_cfg_standard_r_segment_ex_ar_process_inst
      (
      .clk(clk),
      .rst_bar(rst_bar),
      .ar_out_vld(ar_out_vld),
      .ar_out_rdy(ar_out_rdy),
      .ar_out_dat(ar_out_dat),
      .ex_ar_chan_vld(ex_ar_chan_vld),
      .ex_ar_chan_rdy(ex_ar_chan_rdy),
      .ex_ar_chan_dat(ex_ar_chan_dat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    scatter_gather_dma
// ------------------------------------------------------------------


module scatter_gather_dma (
  clk, rst_bar, r_master0_ar_vld, r_master0_ar_rdy, r_master0_ar_dat, r_master0_r_vld,
      r_master0_r_rdy, r_master0_r_dat, w_master0_aw_vld, w_master0_aw_rdy, w_master0_aw_dat,
      w_master0_w_vld, w_master0_w_rdy, w_master0_w_dat, w_master0_b_vld, w_master0_b_rdy,
      w_master0_b_dat, r_slave0_ar_vld, r_slave0_ar_rdy, r_slave0_ar_dat, r_slave0_r_vld,
      r_slave0_r_rdy, r_slave0_r_dat, w_slave0_aw_vld, w_slave0_aw_rdy, w_slave0_aw_dat,
      w_slave0_w_vld, w_slave0_w_rdy, w_slave0_w_dat, w_slave0_b_vld, w_slave0_b_rdy,
      w_slave0_b_dat, dma_done_vld, dma_done_rdy, dma_done_dat
);
  input clk;
  input rst_bar;
  output r_master0_ar_vld;
  input r_master0_ar_rdy;
  output [43:0] r_master0_ar_dat;
  input r_master0_r_vld;
  output r_master0_r_rdy;
  input [70:0] r_master0_r_dat;
  output w_master0_aw_vld;
  input w_master0_aw_rdy;
  output [43:0] w_master0_aw_dat;
  output w_master0_w_vld;
  input w_master0_w_rdy;
  output [72:0] w_master0_w_dat;
  input w_master0_b_vld;
  output w_master0_b_rdy;
  input [5:0] w_master0_b_dat;
  input r_slave0_ar_vld;
  output r_slave0_ar_rdy;
  input [31:0] r_slave0_ar_dat;
  output r_slave0_r_vld;
  input r_slave0_r_rdy;
  output [33:0] r_slave0_r_dat;
  input w_slave0_aw_vld;
  output w_slave0_aw_rdy;
  input [31:0] w_slave0_aw_dat;
  input w_slave0_w_vld;
  output w_slave0_w_rdy;
  input [31:0] w_slave0_w_dat;
  output w_slave0_b_vld;
  input w_slave0_b_rdy;
  output [1:0] w_slave0_b_dat;
  output dma_done_vld;
  input dma_done_rdy;
  output dma_done_dat;


  // Interconnect Declarations
  wire dma_cmd_chan_vld;
  wire dma_cmd_chan_rdy;
  wire [175:0] dma_cmd_chan_dat;
  wire w_segment0_ex_aw_chan_vld;
  wire w_segment0_ex_aw_chan_rdy;
  wire [75:0] w_segment0_ex_aw_chan_dat;
  wire w_segment0_w_chan_vld;
  wire w_segment0_w_chan_rdy;
  wire [72:0] w_segment0_w_chan_dat;
  wire w_segment0_b_chan_vld;
  wire w_segment0_b_chan_rdy;
  wire [5:0] w_segment0_b_chan_dat;
  wire r_segment0_ex_ar_chan_vld;
  wire r_segment0_ex_ar_chan_rdy;
  wire [75:0] r_segment0_ex_ar_chan_dat;


  // Interconnect Declarations for Component Instantiations 
  axi_axi4_segment_axi_cfg_standard_w_segment w_segment0 (
      .clk(clk),
      .rst_bar(rst_bar),
      .aw_out_vld(w_master0_aw_vld),
      .aw_out_rdy(w_master0_aw_rdy),
      .aw_out_dat(w_master0_aw_dat),
      .w_out_vld(w_master0_w_vld),
      .w_out_rdy(w_master0_w_rdy),
      .w_out_dat(w_master0_w_dat),
      .b_in_vld(w_master0_b_vld),
      .b_in_rdy(w_master0_b_rdy),
      .b_in_dat(w_master0_b_dat),
      .ex_aw_chan_vld(w_segment0_ex_aw_chan_vld),
      .ex_aw_chan_rdy(w_segment0_ex_aw_chan_rdy),
      .ex_aw_chan_dat(w_segment0_ex_aw_chan_dat),
      .w_chan_vld(w_segment0_w_chan_vld),
      .w_chan_rdy(w_segment0_w_chan_rdy),
      .w_chan_dat(w_segment0_w_chan_dat),
      .b_chan_vld(w_segment0_b_chan_vld),
      .b_chan_rdy(w_segment0_b_chan_rdy),
      .b_chan_dat(w_segment0_b_chan_dat)
    );
  axi_axi4_segment_axi_cfg_standard_r_segment r_segment0 (
      .clk(clk),
      .rst_bar(rst_bar),
      .ar_out_vld(r_master0_ar_vld),
      .ar_out_rdy(r_master0_ar_rdy),
      .ar_out_dat(r_master0_ar_dat),
      .ex_ar_chan_vld(r_segment0_ex_ar_chan_vld),
      .ex_ar_chan_rdy(r_segment0_ex_ar_chan_rdy),
      .ex_ar_chan_dat(r_segment0_ex_ar_chan_dat)
    );
  scatter_gather_dma_slave_process scatter_gather_dma_slave_process_inst (
      .clk(clk),
      .rst_bar(rst_bar),
      .w_slave0_aw_vld(w_slave0_aw_vld),
      .w_slave0_aw_rdy(w_slave0_aw_rdy),
      .w_slave0_aw_dat(w_slave0_aw_dat),
      .w_slave0_w_vld(w_slave0_w_vld),
      .w_slave0_w_rdy(w_slave0_w_rdy),
      .w_slave0_w_dat(w_slave0_w_dat),
      .w_slave0_b_vld(w_slave0_b_vld),
      .w_slave0_b_rdy(w_slave0_b_rdy),
      .w_slave0_b_dat(w_slave0_b_dat),
      .dma_cmd_chan_vld(dma_cmd_chan_vld),
      .dma_cmd_chan_rdy(dma_cmd_chan_rdy),
      .dma_cmd_chan_dat(dma_cmd_chan_dat)
    );
  scatter_gather_dma_master_process scatter_gather_dma_master_process_inst (
      .clk(clk),
      .rst_bar(rst_bar),
      .r_master0_r_vld(r_master0_r_vld),
      .r_master0_r_rdy(r_master0_r_rdy),
      .r_master0_r_dat(r_master0_r_dat),
      .dma_done_vld(dma_done_vld),
      .dma_done_rdy(dma_done_rdy),
      .dma_done_dat(dma_done_dat),
      .dma_cmd_chan_vld(dma_cmd_chan_vld),
      .dma_cmd_chan_rdy(dma_cmd_chan_rdy),
      .dma_cmd_chan_dat(dma_cmd_chan_dat),
      .w_segment0_ex_aw_chan_vld(w_segment0_ex_aw_chan_vld),
      .w_segment0_ex_aw_chan_rdy(w_segment0_ex_aw_chan_rdy),
      .w_segment0_ex_aw_chan_dat(w_segment0_ex_aw_chan_dat),
      .w_segment0_w_chan_vld(w_segment0_w_chan_vld),
      .w_segment0_w_chan_rdy(w_segment0_w_chan_rdy),
      .w_segment0_w_chan_dat(w_segment0_w_chan_dat),
      .w_segment0_b_chan_vld(w_segment0_b_chan_vld),
      .w_segment0_b_chan_rdy(w_segment0_b_chan_rdy),
      .w_segment0_b_chan_dat(w_segment0_b_chan_dat),
      .r_segment0_ex_ar_chan_vld(r_segment0_ex_ar_chan_vld),
      .r_segment0_ex_ar_chan_rdy(r_segment0_ex_ar_chan_rdy),
      .r_segment0_ex_ar_chan_dat(r_segment0_ex_ar_chan_dat)
    );
  assign r_slave0_ar_rdy = 1'b0;
  assign r_slave0_r_vld = 1'b0;
  assign r_slave0_r_dat = 34'b0000000000000000000000000000000000;
endmodule



