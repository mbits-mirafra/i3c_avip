
import uvm_pkg::*;
import qvip_axi4_bench_test_pkg::*;

module hvl_top;

initial run_test();

endmodule

