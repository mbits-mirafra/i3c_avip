package svdpi;

  import "DPI-C" context function chandle svGetScopeFromName ( input string path );
  import "DPI-C" context function string svGetNameFromScope( input chandle scope );

endpackage
