//
// File: hvl_scatter_gather_dma_qvip.sv
//
// Generated from Mentor VIP Configurator (20201007)
// Generated using Mentor VIP Library ( 2020.4 : 10/16/2020:13:17 )
//
module hvl_scatter_gather_dma_qvip;
    import uvm_pkg::*;
    
    `include "test_packages.svh"
    
    initial
    begin
        run_test();
    end

endmodule: hvl_scatter_gather_dma_qvip
