//
// File: hvl_axi4_2x2_fabric_qvip.sv
//
// Generated from Mentor VIP Configurator (20191003)
// Generated using Mentor VIP Library ( 2019.4 : 10/16/2019:13:47 )
//
module hvl_axi4_2x2_fabric_qvip;
    import uvm_pkg::*;
    
    `include "test_packages.svh"
    
    initial
    begin
        run_test();
    end

endmodule: hvl_axi4_2x2_fabric_qvip
