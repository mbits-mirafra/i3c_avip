//----------------------------------------------------------------------
// Created with uvmf_gen version 2019.4_1
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef enum {SPI_SLAVE_READ, SPI_SLAVE_WRITE} spi_op_t;
typedef enum {MOSI, MISO, TO_SPI, FROM_SPI} spi_dir_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

