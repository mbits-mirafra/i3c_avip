//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This environment contains all agents, predictors and
// scoreboards required for the block level design.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

class env_environment  extends uvmf_environment_base #(
    .CONFIG_T( env_env_configuration 
  ));
  `uvm_component_utils( env_environment )





  typedef i3c_m_agent  m_agent_t;
  m_agent_t m_agent;

  typedef i3c_s_agent  s_agent_t;
  s_agent_t s_agent;




  typedef i3c_scoreboard #(
                .CONFIG_T(CONFIG_T)
                ) i3c_sb_t;
  i3c_sb_t i3c_sb;




  typedef uvmf_virtual_sequencer_base #(.CONFIG_T(env_env_configuration)) env_vsqr_t;
  env_vsqr_t vsqr;

  // pragma uvmf custom class_item_additional begin
  // pragma uvmf custom class_item_additional end
 
// ****************************************************************************
// FUNCTION : new()
// This function is the standard SystemVerilog constructor.
//
  function new( string name = "", uvm_component parent = null );
    super.new( name, parent );
  endfunction

// ****************************************************************************
// FUNCTION: build_phase()
// This function builds all components within this environment.
//
  virtual function void build_phase(uvm_phase phase);
// pragma uvmf custom build_phase_pre_super begin
// pragma uvmf custom build_phase_pre_super end
    super.build_phase(phase);
    m_agent = m_agent_t::type_id::create("m_agent",this);
    m_agent.set_config(configuration.m_agent_config);
    s_agent = s_agent_t::type_id::create("s_agent",this);
    s_agent.set_config(configuration.s_agent_config);
    i3c_sb = i3c_sb_t::type_id::create("i3c_sb",this);
    i3c_sb.configuration = configuration;

    vsqr = env_vsqr_t::type_id::create("vsqr", this);
    vsqr.set_config(configuration);
    configuration.set_vsqr(vsqr);

    // pragma uvmf custom build_phase begin
    // pragma uvmf custom build_phase end
  endfunction

// ****************************************************************************
// FUNCTION: connect_phase()
// This function makes all connections within this environment.  Connections
// typically inclue agent to predictor, predictor to scoreboard and scoreboard
// to agent.
//
  virtual function void connect_phase(uvm_phase phase);
// pragma uvmf custom connect_phase_pre_super begin
// pragma uvmf custom connect_phase_pre_super end
    super.connect_phase(phase);
    m_agent.monitored_ap.connect(i3c_sb.m_sb_ep);
    s_agent.monitored_ap.connect(i3c_sb.s_sb_ep);
    // pragma uvmf custom reg_model_connect_phase begin
    // pragma uvmf custom reg_model_connect_phase end
  endfunction

// ****************************************************************************
// FUNCTION: end_of_simulation_phase()
// This function is executed just prior to executing run_phase.  This function
// was added to the environment to sample environment configuration settings
// just before the simulation exits time 0.  The configuration structure is 
// randomized in the build phase before the environment structure is constructed.
// Configuration variables can be customized after randomization in the build_phase
// of the extended test.
// If a sequence modifies values in the configuration structure then the sequence is
// responsible for sampling the covergroup in the configuration if required.
//
  virtual function void start_of_simulation_phase(uvm_phase phase);
     configuration.env_configuration_cg.sample();
  endfunction

endclass

// pragma uvmf custom external begin
// pragma uvmf custom external end

