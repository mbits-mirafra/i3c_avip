`ifndef I3C_CONTROLLER_READOPERATIONWITHRANDOMDATATRANSFERWIDTH_SEQ_INCLUDED_
`define I3C_CONTROLLER_READOPERATIONWITHRANDOMDATATRANSFERWIDTH_SEQ_INCLUDED_

class i3c_controller_readOperationWithRandomDataTransferWidth_seq extends i3c_controller_base_seq;
  `uvm_object_utils(i3c_controller_readOperationWithRandomDataTransferWidth_seq)

  extern function new(string name = "i3c_controller_readOperationWithRandomDataTransferWidth_seq");
  extern task body();
endclass : i3c_controller_readOperationWithRandomDataTransferWidth_seq

function i3c_controller_readOperationWithRandomDataTransferWidth_seq::new(string name = "i3c_controller_readOperationWithRandomDataTransferWidth_seq");
  super.new(name);
endfunction : new


task i3c_controller_readOperationWithRandomDataTransferWidth_seq::body();
  super.body();

  req = i3c_controller_tx::type_id::create("req"); 

  start_item(req);
    if(!req.randomize() with {operation == READ;
                              targetAddress == 7'b1010101;}) begin
      `uvm_error(get_type_name(), "Randomization failed")
    end
  
    req.print();
  finish_item(req);

endtask:body
  
`endif


