`ifndef I3C_CONTROLLER_BASE_SEQ_INCLUDED_
`define I3C_CONTROLLER_BASE_SEQ_INCLUDED_

class i3c_controller_base_seq extends uvm_sequence #(i3c_controller_tx);
  `uvm_object_utils(i3c_controller_base_seq)

  // GopalS:  `uvm_declare_p_sequencer(i3c_controller_sequencer) 

  extern function new(string name = "i3c_controller_base_seq");
  extern virtual task body();
endclass : i3c_controller_base_seq


function i3c_controller_base_seq::new(string name = "i3c_controller_base_seq");
  super.new(name);
endfunction : new

task i3c_controller_base_seq::body();
//super.body();
//dynamic casting of p_sequencer and m_sequencer
// GopalS:    if(!$cast(p_sequencer,m_sequencer))begin
// GopalS:      `uvm_error(get_full_name(),"Virtual sequencer pointer cast failed")
// GopalS:    end
            
endtask:body

`endif
