//----------------------------------------------------------------------
// Created with uvmf_gen version 2019.4_1
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This file contains macros used with the gpio package.
//   These macros include packed struct definitions.  These structs are
//   used to pass data between classes, hvl, and BFM's, hdl.  Use of 
//   structs are more efficient and simpler to modify.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_struct
//      and from_struct methods defined in the macros below that are used in  
//      the gpio_configuration class.
//
  `define gpio_CONFIGURATION_STRUCT \
typedef struct packed  { \
     uvmf_active_passive_t active_passive; \
     uvmf_initiator_responder_t initiator_responder; \
     } gpio_configuration_s;

  `define gpio_CONFIGURATION_TO_STRUCT_FUNCTION \
  virtual function gpio_configuration_s to_struct();\
    gpio_configuration_struct = \
       {\
       this.active_passive,\
       this.initiator_responder\
       };\
    return ( gpio_configuration_struct );\
  endfunction

  `define gpio_CONFIGURATION_FROM_STRUCT_FUNCTION \
  virtual function void from_struct(gpio_configuration_s gpio_configuration_struct);\
      {\
      this.active_passive,\
      this.initiator_responder  \
      } = gpio_configuration_struct;\
  endfunction

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_monitor_struct
//      and from_monitor_struct methods of the gpio_transaction class.
//
  `define gpio_MONITOR_STRUCT typedef struct packed  { \
  gpio_op_t op ; \
  logic [READ_PORT_WIDTH-1:0] read_port ; \
  logic [WRITE_PORT_WIDTH-1:0] write_port ; \
     } gpio_monitor_s;

  `define gpio_TO_MONITOR_STRUCT_FUNCTION \
  virtual function gpio_monitor_s to_monitor_struct();\
    gpio_monitor_struct = \
            { \
            this.op , \
            this.read_port , \
            this.write_port  \
            };\
    return ( gpio_monitor_struct);\
  endfunction\

  `define gpio_FROM_MONITOR_STRUCT_FUNCTION \
  virtual function void from_monitor_struct(gpio_monitor_s gpio_monitor_struct);\
            {\
            this.op , \
            this.read_port , \
            this.write_port  \
            } = gpio_monitor_struct;\
  endfunction

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_initiator_struct
//      and from_initiator_struct methods of the gpio_transaction class.
//      Also update the comments in the driver BFM.
//
  `define gpio_INITIATOR_STRUCT typedef struct packed  { \
  gpio_op_t op ; \
  logic [READ_PORT_WIDTH-1:0] read_port ; \
  logic [WRITE_PORT_WIDTH-1:0] write_port ; \
     } gpio_initiator_s;

  `define gpio_TO_INITIATOR_STRUCT_FUNCTION \
  virtual function gpio_initiator_s to_initiator_struct();\
    gpio_initiator_struct = \
           {\
           this.op , \
           this.read_port , \
           this.write_port  \
           };\
    return ( gpio_initiator_struct);\
  endfunction

  `define gpio_FROM_INITIATOR_STRUCT_FUNCTION \
  virtual function void from_initiator_struct(gpio_initiator_s gpio_initiator_struct);\
           {\
           this.op , \
           this.read_port , \
           this.write_port  \
           } = gpio_initiator_struct;\
  endfunction

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_responder_struct
//      and from_responder_struct methods of the gpio_transaction class.
//      Also update the comments in the driver BFM.
//
  `define gpio_RESPONDER_STRUCT typedef struct packed  { \
  gpio_op_t op ; \
  logic [READ_PORT_WIDTH-1:0] read_port ; \
  logic [WRITE_PORT_WIDTH-1:0] write_port ; \
     } gpio_responder_s;

  `define gpio_TO_RESPONDER_STRUCT_FUNCTION \
  virtual function gpio_responder_s to_responder_struct();\
    gpio_responder_struct = \
           {\
           this.op , \
           this.read_port , \
           this.write_port  \
           };\
    return ( gpio_responder_struct);\
  endfunction

  `define gpio_FROM_RESPONDER_STRUCT_FUNCTION \
  virtual function void from_responder_struct(gpio_responder_s gpio_responder_struct);\
           {\
           this.op , \
           this.read_port , \
           this.write_port  \
           } = gpio_responder_struct;\
  endfunction
// pragma uvmf custom additional begin
// pragma uvmf custom additional end
