//
// File: test_packages.svh
//
// Generated from Mentor VIP Configurator (20201007)
// Generated using Mentor VIP Library ( 2020.4 : 10/16/2020:13:17 )
//

import scatter_gather_dma_qvip_pkg::*;

// Add other packages here as required
