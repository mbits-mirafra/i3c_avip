import "DPI-C" context function void trigger_hvl_event(int unsigned ret_val = 0);
import "DPI-C" context function void trigger_numbered_hvl_event(int unsigned event_num, int unsigned ret_val = 0);
