//
// File: scatter_gather_dma_qvip_pkg.sv
//
// Generated from Mentor VIP Configurator (20201007)
// Generated using Mentor VIP Library ( 2020.4 : 10/16/2020:13:17 )
//
package scatter_gather_dma_qvip_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    
    import addr_map_pkg::*;
    
    import scatter_gather_dma_qvip_params_pkg::*;
    import mvc_pkg::*;
    import mgc_axi4_v1_0_pkg::*;
    
    `include "scatter_gather_dma_qvip_env_config.svh"
    `include "scatter_gather_dma_qvip_env.svh"
    `include "scatter_gather_dma_qvip_vseq_base.svh"
    `include "scatter_gather_dma_qvip_test_base.svh"
endpackage: scatter_gather_dma_qvip_pkg
