//----------------------------------------------------------------------
//   Copyright 2013 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//                   Mentor Graphics Inc
//----------------------------------------------------------------------
// Project         : APB3
// Unit            : APB3 Memory Slave Module
// File            : apb3_memory_slave_module.svh
//----------------------------------------------------------------------
// Creation Date   : 07.25.2013
//----------------------------------------------------------------------
// Description: This module implements a memory slave for the apb3 bus.
//    It is a self contained module that can be attached to an mgc_apb3
//    interface as an rtl slave.
//
//----------------------------------------------------------------------
//

`include "uvm_macros.svh"

module apb3_memory_slave_module(PCLK, PRESETn, PADDR, PSEL, PENABLE, PWRITE, PWDATA, PRDATA, PREADY, PSLVERR);
  import uvm_pkg::*;
  import mvc_pkg::*;
  import mgc_apb3_v1_0_pkg::*;

  parameter ADDRESS_WIDTH = 32;
  parameter WDATA_WIDTH   = 32;
  parameter RDATA_WIDTH   = 32;
  parameter AGENT_NAME = "";

  // system signals
  input PCLK   ;
  input PRESETn;

  // Slave input signals
  input [ADDRESS_WIDTH-1:0] PADDR;
  input                     PSEL;
  input                     PENABLE;
  input                     PWRITE;
  input [WDATA_WIDTH-1:0]   PWDATA;

  // Slave output signals
  output [RDATA_WIDTH-1:0]  PRDATA;
  output                    PREADY;
  output                    PSLVERR;

 
  string agent_name = (AGENT_NAME == "")? $psprintf("%m") : 
  `ifdef MODEL_TECH 
    AGENT_NAME;
  `else
    $psprintf("%s",AGENT_NAME);
  `endif

  mgc_apb3 #(1, ADDRESS_WIDTH, WDATA_WIDTH, RDATA_WIDTH) apb3_if(PCLK, PRESETn);

  // Signals driven by slave
  assign PREADY  = (PSEL)? apb3_if.PREADY  : 'bz;
  assign PRDATA  = (PSEL)? apb3_if.PRDATA  : 'bz;
  assign PSLVERR = (PSEL)? apb3_if.PSLVERR : 'bz;

  // Signals driven by master
  assign apb3_if.PADDR   = PADDR;
  assign apb3_if.PSEL     = PSEL;
  assign apb3_if.PENABLE  = PENABLE;
  assign apb3_if.PWRITE   = PWRITE;
  assign apb3_if.PWDATA   = PWDATA;

`ifdef APB3_QVL_MONITOR
  qvl_amba3_apb_monitor #(
                          .ADD_BUS_WIDTH(ADDRESS_WIDTH), 
                          .DATA_BUS_WIDTH((WDATA_WIDTH > RDATA_WIDTH)? RDATA_WIDTH : WDATA_WIDTH)
                         )
                 slave_qvl(
                           .pclk(apb3_if.PCLK), 
                           .presetn(apb3_if.PRESETn), 
                           .paddr(apb3_if.PADDR), 
                           .pselx(apb3_if.PSEL), 
                           .penable(apb3_if.PENABLE),
                           .pwrite(apb3_if.PWRITE), 
                           .pwdata(apb3_if.PWDATA), 
                           .prdata(apb3_if.PRDATA),
                           .pready(apb3_if.PREADY),
                           .pslverr(apb3_if.PSLVERR)
                          );
`endif

  initial begin
    uvm_object o;
    uvm_root top;
    mvc_env_config c;
    apb3_vip_config #(1 , ADDRESS_WIDTH , WDATA_WIDTH , RDATA_WIDTH) slave_config;

    top = uvm_root::get();

    if(!uvm_config_db #( uvm_object )::get( top , "" , s_top_level_config_id , o))
    begin
      c = new();
    end
    else
    begin
      if ( !$cast(c , o) )  
        `uvm_fatal("CONFIG_EROR" ,
                           $psprintf( "config with id must be of type top_level_config") );
    end

    slave_config = new();
    slave_config.m_bfm = apb3_if;

    // Master is RTL, slave is TLM
    slave_config.m_bfm.apb3_set_host_abstraction_level(1, 0);
    slave_config.m_bfm.apb3_set_slave_abstraction_level(0, 1);
     
    // Clocks and resets generated by RTL;
    slave_config.m_bfm.apb3_set_clk_contr_abstraction_level(1, 0);
    slave_config.m_bfm.apb3_set_rst_contr_abstraction_level(1, 0);

    // Add Memory slave functionality
    slave_config.set_default_sequence(apb3_transaction_memory_sequence #(1, ADDRESS_WIDTH, WDATA_WIDTH, RDATA_WIDTH)::get_type(), 1); 

    apb3_if._initialized();

    c.add_child_config(agent_name, slave_config);
    uvm_config_db #( uvm_object )::set( null , "*" , s_top_level_config_id , c );
  end

endmodule

           

